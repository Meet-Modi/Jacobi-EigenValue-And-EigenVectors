`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:12:13 11/09/2018 
// Design Name: 
// Module Name:    Matrix_Multiply_32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Matrix_Multiply_32(select_line_in, A_wire, B_wire,index_A, index_B, clk, reset, out, out_address, select_line_out, write_data);
	output reg [1023:0] out;
	output reg [4:0] out_address;
	output reg select_line_out, write_data;
	input select_line_in;
	input clk, reset; 
	input [1023:0] A_wire, B_wire;
	input [4:0] index_A, index_B;
	reg [31:0] A [0:31][0:31];
	reg [31:0] B [0:31][0:31];
	reg [31:0] C [0:31][0:31];
	wire [5:0] counter;
	reg [5:0] counter_reg;
	reg loaded_flag;
	reg [5:0] i;
	reg [4:0] address_reg;
	wire [4:0] address;
	
	wire [31:0] mul0, mul1, mul2, mul3, mul4, mul5, mul6, mul7, mul8, mul9, mul10, mul11, mul12, mul13, mul14, mul15, mul16, mul17, mul18, mul19, mul20, mul21, mul22, mul23, mul24, mul25, mul26, mul27, mul28, mul29, mul30, mul31 ;
	wire [31:0] mul32, mul33, mul34, mul35, mul36, mul37, mul38, mul39, mul40, mul41, mul42, mul43, mul44, mul45, mul46, mul47, mul48, mul49, mul50, mul51, mul52, mul53, mul54, mul55, mul56, mul57, mul58, mul59, mul60, mul61, mul62, mul63 ;
	wire [31:0] mul64, mul65, mul66, mul67, mul68, mul69, mul70, mul71, mul72, mul73, mul74, mul75, mul76, mul77, mul78, mul79, mul80, mul81, mul82, mul83, mul84, mul85, mul86, mul87, mul88, mul89, mul90, mul91, mul92, mul93, mul94, mul95 ;
	wire [31:0] mul96, mul97, mul98, mul99, mul100, mul101, mul102, mul103, mul104, mul105, mul106, mul107, mul108, mul109, mul110, mul111, mul112, mul113, mul114, mul115, mul116, mul117, mul118, mul119, mul120, mul121, mul122, mul123, mul124, mul125, mul126, mul127 ;
	wire [31:0] mul128, mul129, mul130, mul131, mul132, mul133, mul134, mul135, mul136, mul137, mul138, mul139, mul140, mul141, mul142, mul143, mul144, mul145, mul146, mul147, mul148, mul149, mul150, mul151, mul152, mul153, mul154, mul155, mul156, mul157, mul158, mul159 ;
	wire [31:0] mul160, mul161, mul162, mul163, mul164, mul165, mul166, mul167, mul168, mul169, mul170, mul171, mul172, mul173, mul174, mul175, mul176, mul177, mul178, mul179, mul180, mul181, mul182, mul183, mul184, mul185, mul186, mul187, mul188, mul189, mul190, mul191 ;
	wire [31:0] mul192, mul193, mul194, mul195, mul196, mul197, mul198, mul199, mul200, mul201, mul202, mul203, mul204, mul205, mul206, mul207, mul208, mul209, mul210, mul211, mul212, mul213, mul214, mul215, mul216, mul217, mul218, mul219, mul220, mul221, mul222, mul223 ;
	wire [31:0] mul224, mul225, mul226, mul227, mul228, mul229, mul230, mul231, mul232, mul233, mul234, mul235, mul236, mul237, mul238, mul239, mul240, mul241, mul242, mul243, mul244, mul245, mul246, mul247, mul248, mul249, mul250, mul251, mul252, mul253, mul254, mul255 ;
	wire [31:0] mul256, mul257, mul258, mul259, mul260, mul261, mul262, mul263, mul264, mul265, mul266, mul267, mul268, mul269, mul270, mul271, mul272, mul273, mul274, mul275, mul276, mul277, mul278, mul279, mul280, mul281, mul282, mul283, mul284, mul285, mul286, mul287 ;
	wire [31:0] mul288, mul289, mul290, mul291, mul292, mul293, mul294, mul295, mul296, mul297, mul298, mul299, mul300, mul301, mul302, mul303, mul304, mul305, mul306, mul307, mul308, mul309, mul310, mul311, mul312, mul313, mul314, mul315, mul316, mul317, mul318, mul319 ;
	wire [31:0] mul320, mul321, mul322, mul323, mul324, mul325, mul326, mul327, mul328, mul329, mul330, mul331, mul332, mul333, mul334, mul335, mul336, mul337, mul338, mul339, mul340, mul341, mul342, mul343, mul344, mul345, mul346, mul347, mul348, mul349, mul350, mul351 ;
	wire [31:0] mul352, mul353, mul354, mul355, mul356, mul357, mul358, mul359, mul360, mul361, mul362, mul363, mul364, mul365, mul366, mul367, mul368, mul369, mul370, mul371, mul372, mul373, mul374, mul375, mul376, mul377, mul378, mul379, mul380, mul381, mul382, mul383 ;
	wire [31:0] mul384, mul385, mul386, mul387, mul388, mul389, mul390, mul391, mul392, mul393, mul394, mul395, mul396, mul397, mul398, mul399, mul400, mul401, mul402, mul403, mul404, mul405, mul406, mul407, mul408, mul409, mul410, mul411, mul412, mul413, mul414, mul415 ;
	wire [31:0] mul416, mul417, mul418, mul419, mul420, mul421, mul422, mul423, mul424, mul425, mul426, mul427, mul428, mul429, mul430, mul431, mul432, mul433, mul434, mul435, mul436, mul437, mul438, mul439, mul440, mul441, mul442, mul443, mul444, mul445, mul446, mul447 ;
	wire [31:0] mul448, mul449, mul450, mul451, mul452, mul453, mul454, mul455, mul456, mul457, mul458, mul459, mul460, mul461, mul462, mul463, mul464, mul465, mul466, mul467, mul468, mul469, mul470, mul471, mul472, mul473, mul474, mul475, mul476, mul477, mul478, mul479 ;
	wire [31:0] mul480, mul481, mul482, mul483, mul484, mul485, mul486, mul487, mul488, mul489, mul490, mul491, mul492, mul493, mul494, mul495, mul496, mul497, mul498, mul499, mul500, mul501, mul502, mul503, mul504, mul505, mul506, mul507, mul508, mul509, mul510, mul511 ;
	wire [31:0] mul512, mul513, mul514, mul515, mul516, mul517, mul518, mul519, mul520, mul521, mul522, mul523, mul524, mul525, mul526, mul527, mul528, mul529, mul530, mul531, mul532, mul533, mul534, mul535, mul536, mul537, mul538, mul539, mul540, mul541, mul542, mul543 ;
	wire [31:0] mul544, mul545, mul546, mul547, mul548, mul549, mul550, mul551, mul552, mul553, mul554, mul555, mul556, mul557, mul558, mul559, mul560, mul561, mul562, mul563, mul564, mul565, mul566, mul567, mul568, mul569, mul570, mul571, mul572, mul573, mul574, mul575 ;
	wire [31:0] mul576, mul577, mul578, mul579, mul580, mul581, mul582, mul583, mul584, mul585, mul586, mul587, mul588, mul589, mul590, mul591, mul592, mul593, mul594, mul595, mul596, mul597, mul598, mul599, mul600, mul601, mul602, mul603, mul604, mul605, mul606, mul607 ;
	wire [31:0] mul608, mul609, mul610, mul611, mul612, mul613, mul614, mul615, mul616, mul617, mul618, mul619, mul620, mul621, mul622, mul623, mul624, mul625, mul626, mul627, mul628, mul629, mul630, mul631, mul632, mul633, mul634, mul635, mul636, mul637, mul638, mul639 ;
	wire [31:0] mul640, mul641, mul642, mul643, mul644, mul645, mul646, mul647, mul648, mul649, mul650, mul651, mul652, mul653, mul654, mul655, mul656, mul657, mul658, mul659, mul660, mul661, mul662, mul663, mul664, mul665, mul666, mul667, mul668, mul669, mul670, mul671 ;
	wire [31:0] mul672, mul673, mul674, mul675, mul676, mul677, mul678, mul679, mul680, mul681, mul682, mul683, mul684, mul685, mul686, mul687, mul688, mul689, mul690, mul691, mul692, mul693, mul694, mul695, mul696, mul697, mul698, mul699, mul700, mul701, mul702, mul703 ;
	wire [31:0] mul704, mul705, mul706, mul707, mul708, mul709, mul710, mul711, mul712, mul713, mul714, mul715, mul716, mul717, mul718, mul719, mul720, mul721, mul722, mul723, mul724, mul725, mul726, mul727, mul728, mul729, mul730, mul731, mul732, mul733, mul734, mul735 ;
	wire [31:0] mul736, mul737, mul738, mul739, mul740, mul741, mul742, mul743, mul744, mul745, mul746, mul747, mul748, mul749, mul750, mul751, mul752, mul753, mul754, mul755, mul756, mul757, mul758, mul759, mul760, mul761, mul762, mul763, mul764, mul765, mul766, mul767 ;
	wire [31:0] mul768, mul769, mul770, mul771, mul772, mul773, mul774, mul775, mul776, mul777, mul778, mul779, mul780, mul781, mul782, mul783, mul784, mul785, mul786, mul787, mul788, mul789, mul790, mul791, mul792, mul793, mul794, mul795, mul796, mul797, mul798, mul799 ;
	wire [31:0] mul800, mul801, mul802, mul803, mul804, mul805, mul806, mul807, mul808, mul809, mul810, mul811, mul812, mul813, mul814, mul815, mul816, mul817, mul818, mul819, mul820, mul821, mul822, mul823, mul824, mul825, mul826, mul827, mul828, mul829, mul830, mul831 ;
	wire [31:0] mul832, mul833, mul834, mul835, mul836, mul837, mul838, mul839, mul840, mul841, mul842, mul843, mul844, mul845, mul846, mul847, mul848, mul849, mul850, mul851, mul852, mul853, mul854, mul855, mul856, mul857, mul858, mul859, mul860, mul861, mul862, mul863 ;
	wire [31:0] mul864, mul865, mul866, mul867, mul868, mul869, mul870, mul871, mul872, mul873, mul874, mul875, mul876, mul877, mul878, mul879, mul880, mul881, mul882, mul883, mul884, mul885, mul886, mul887, mul888, mul889, mul890, mul891, mul892, mul893, mul894, mul895 ;
	wire [31:0] mul896, mul897, mul898, mul899, mul900, mul901, mul902, mul903, mul904, mul905, mul906, mul907, mul908, mul909, mul910, mul911, mul912, mul913, mul914, mul915, mul916, mul917, mul918, mul919, mul920, mul921, mul922, mul923, mul924, mul925, mul926, mul927 ;
	wire [31:0] mul928, mul929, mul930, mul931, mul932, mul933, mul934, mul935, mul936, mul937, mul938, mul939, mul940, mul941, mul942, mul943, mul944, mul945, mul946, mul947, mul948, mul949, mul950, mul951, mul952, mul953, mul954, mul955, mul956, mul957, mul958, mul959 ;
	wire [31:0] mul960, mul961, mul962, mul963, mul964, mul965, mul966, mul967, mul968, mul969, mul970, mul971, mul972, mul973, mul974, mul975, mul976, mul977, mul978, mul979, mul980, mul981, mul982, mul983, mul984, mul985, mul986, mul987, mul988, mul989, mul990, mul991 ;
	wire [31:0] mul992, mul993, mul994, mul995, mul996, mul997, mul998, mul999, mul1000, mul1001, mul1002, mul1003, mul1004, mul1005, mul1006, mul1007, mul1008, mul1009, mul1010, mul1011, mul1012, mul1013, mul1014, mul1015, mul1016, mul1017, mul1018, mul1019, mul1020, mul1021, mul1022, mul1023 ;
	wire [31:0] s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43, s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57, s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71, s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85, s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99, s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111, s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123, s124, s125, s126, s127, s128, s129, s130, s131, s132, s133, s134, s135, s136, s137, s138, s139, s140, s141, s142, s143, s144, s145, s146, s147, s148, s149, s150, s151, s152, s153, s154, s155, s156, s157, s158, s159, s160, s161, s162, s163, s164, s165, s166, s167, s168, s169, s170, s171, s172, s173, s174, s175, s176, s177, s178, s179, s180, s181, s182, s183, s184, s185, s186, s187, s188, s189, s190, s191, s192, s193, s194, s195, s196, s197, s198, s199, s200, s201, s202, s203, s204, s205, s206, s207, s208, s209, s210, s211, s212, s213, s214, s215, s216, s217, s218, s219, s220, s221, s222, s223, s224, s225, s226, s227, s228, s229, s230, s231, s232, s233, s234, s235, s236, s237, s238, s239, s240, s241, s242, s243, s244, s245, s246, s247, s248, s249, s250, s251, s252, s253, s254, s255, s256, s257, s258, s259, s260, s261, s262, s263, s264, s265, s266, s267, s268, s269, s270, s271, s272, s273, s274, s275, s276, s277, s278, s279, s280, s281, s282, s283, s284, s285, s286, s287, s288, s289, s290, s291, s292, s293, s294, s295, s296, s297, s298, s299, s300, s301, s302, s303, s304, s305, s306, s307, s308, s309, s310, s311, s312, s313, s314, s315, s316, s317, s318, s319, s320, s321, s322, s323, s324, s325, s326, s327, s328, s329, s330, s331, s332, s333, s334, s335, s336, s337, s338, s339, s340, s341, s342, s343, s344, s345, s346, s347, s348, s349, s350, s351, s352, s353, s354, s355, s356, s357, s358, s359, s360, s361, s362, s363, s364, s365, s366, s367, s368, s369, s370, s371, s372, s373, s374, s375, s376, s377, s378, s379, s380, s381, s382, s383, s384, s385, s386, s387, s388, s389, s390, s391, s392, s393, s394, s395, s396, s397, s398, s399, s400, s401, s402, s403, s404, s405, s406, s407, s408, s409, s410, s411, s412, s413, s414, s415, s416, s417, s418, s419, s420, s421, s422, s423, s424, s425, s426, s427, s428, s429, s430, s431, s432, s433, s434, s435, s436, s437, s438, s439, s440, s441, s442, s443, s444, s445, s446, s447, s448, s449, s450, s451, s452, s453, s454, s455, s456, s457, s458, s459, s460, s461, s462, s463, s464, s465, s466, s467, s468, s469, s470, s471, s472, s473, s474, s475, s476, s477, s478, s479, s480, s481, s482, s483, s484, s485, s486, s487, s488, s489, s490, s491, s492, s493, s494, s495, s496, s497, s498, s499, s500, s501, s502, s503, s504, s505, s506, s507, s508, s509, s510, s511, s512, s513, s514, s515, s516, s517, s518, s519, s520, s521, s522, s523, s524, s525, s526, s527, s528, s529, s530, s531, s532, s533, s534, s535, s536, s537, s538, s539, s540, s541, s542, s543, s544, s545, s546, s547, s548, s549, s550, s551, s552, s553, s554, s555, s556, s557, s558, s559, s560, s561, s562, s563, s564, s565, s566, s567, s568, s569, s570, s571, s572, s573, s574, s575, s576, s577, s578, s579, s580, s581, s582, s583, s584, s585, s586, s587, s588, s589, s590, s591, s592, s593, s594, s595, s596, s597, s598, s599, s600, s601, s602, s603, s604, s605, s606, s607, s608, s609, s610, s611, s612, s613, s614, s615, s616, s617, s618, s619, s620, s621, s622, s623, s624, s625, s626, s627, s628, s629, s630, s631, s632, s633, s634, s635, s636, s637, s638, s639, s640, s641, s642, s643, s644, s645, s646, s647, s648, s649, s650, s651, s652, s653, s654, s655, s656, s657, s658, s659, s660, s661, s662, s663, s664, s665, s666, s667, s668, s669, s670, s671, s672, s673, s674, s675, s676, s677, s678, s679, s680, s681, s682, s683, s684, s685, s686, s687, s688, s689, s690, s691, s692, s693, s694, s695, s696, s697, s698, s699, s700, s701, s702, s703, s704, s705, s706, s707, s708, s709, s710, s711, s712, s713, s714, s715, s716, s717, s718, s719, s720, s721, s722, s723, s724, s725, s726, s727, s728, s729, s730, s731, s732, s733, s734, s735, s736, s737, s738, s739, s740, s741, s742, s743, s744, s745, s746, s747, s748, s749, s750, s751, s752, s753, s754, s755, s756, s757, s758, s759, s760, s761, s762, s763, s764, s765, s766, s767, s768, s769, s770, s771, s772, s773, s774, s775, s776, s777, s778, s779, s780, s781, s782, s783, s784, s785, s786, s787, s788, s789, s790, s791, s792, s793, s794, s795, s796, s797, s798, s799, s800, s801, s802, s803, s804, s805, s806, s807, s808, s809, s810, s811, s812, s813, s814, s815, s816, s817, s818, s819, s820, s821, s822, s823, s824, s825, s826, s827, s828, s829, s830, s831, s832, s833, s834, s835, s836, s837, s838, s839, s840, s841, s842, s843, s844, s845, s846, s847, s848, s849, s850, s851, s852, s853, s854, s855, s856, s857, s858, s859, s860, s861, s862, s863, s864, s865, s866, s867, s868, s869, s870, s871, s872, s873, s874, s875, s876, s877, s878, s879, s880, s881, s882, s883, s884, s885, s886, s887, s888, s889, s890, s891, s892, s893, s894, s895, s896, s897, s898, s899, s900, s901, s902, s903, s904, s905, s906, s907, s908, s909, s910, s911, s912, s913, s914, s915, s916, s917, s918, s919, s920, s921, s922, s923, s924, s925, s926, s927, s928, s929, s930, s931, s932, s933, s934, s935, s936, s937, s938, s939, s940, s941, s942, s943, s944, s945, s946, s947, s948, s949, s950, s951, s952, s953, s954, s955, s956, s957, s958, s959, s960, s961, s962, s963, s964, s965, s966, s967, s968, s969, s970, s971, s972, s973, s974, s975, s976, s977, s978, s979, s980, s981, s982, s983, s984, s985, s986, s987, s988, s989, s990, s991;

	multiplier m0(A[address][0],B[0][0],mul0);   multiplier m1(A[address][1],B[1][0],mul1);   multiplier m2(A[address][2],B[2][0],mul2);   multiplier m3(A[address][3],B[3][0],mul3);   multiplier m4(A[address][4],B[4][0],mul4);   multiplier m5(A[address][5],B[5][0],mul5);   multiplier m6(A[address][6],B[6][0],mul6);   multiplier m7(A[address][7],B[7][0],mul7);   multiplier m8(A[address][8],B[8][0],mul8);   multiplier m9(A[address][9],B[9][0],mul9);   multiplier m10(A[address][10],B[10][0],mul10);   multiplier m11(A[address][11],B[11][0],mul11);   multiplier m12(A[address][12],B[12][0],mul12);   multiplier m13(A[address][13],B[13][0],mul13);   multiplier m14(A[address][14],B[14][0],mul14);   multiplier m15(A[address][15],B[15][0],mul15);   multiplier m16(A[address][16],B[16][0],mul16);   multiplier m17(A[address][17],B[17][0],mul17);   multiplier m18(A[address][18],B[18][0],mul18);   multiplier m19(A[address][19],B[19][0],mul19);   multiplier m20(A[address][20],B[20][0],mul20);   multiplier m21(A[address][21],B[21][0],mul21);   multiplier m22(A[address][22],B[22][0],mul22);   multiplier m23(A[address][23],B[23][0],mul23);   multiplier m24(A[address][24],B[24][0],mul24);   multiplier m25(A[address][25],B[25][0],mul25);   multiplier m26(A[address][26],B[26][0],mul26);   multiplier m27(A[address][27],B[27][0],mul27);   multiplier m28(A[address][28],B[28][0],mul28);   multiplier m29(A[address][29],B[29][0],mul29);   multiplier m30(A[address][30],B[30][0],mul30);   multiplier m31(A[address][31],B[31][0],mul31);   
	multiplier m32(A[address][0],B[0][1],mul32);   multiplier m33(A[address][1],B[1][1],mul33);   multiplier m34(A[address][2],B[2][1],mul34);   multiplier m35(A[address][3],B[3][1],mul35);   multiplier m36(A[address][4],B[4][1],mul36);   multiplier m37(A[address][5],B[5][1],mul37);   multiplier m38(A[address][6],B[6][1],mul38);   multiplier m39(A[address][7],B[7][1],mul39);   multiplier m40(A[address][8],B[8][1],mul40);   multiplier m41(A[address][9],B[9][1],mul41);   multiplier m42(A[address][10],B[10][1],mul42);   multiplier m43(A[address][11],B[11][1],mul43);   multiplier m44(A[address][12],B[12][1],mul44);   multiplier m45(A[address][13],B[13][1],mul45);   multiplier m46(A[address][14],B[14][1],mul46);   multiplier m47(A[address][15],B[15][1],mul47);   multiplier m48(A[address][16],B[16][1],mul48);   multiplier m49(A[address][17],B[17][1],mul49);   multiplier m50(A[address][18],B[18][1],mul50);   multiplier m51(A[address][19],B[19][1],mul51);   multiplier m52(A[address][20],B[20][1],mul52);   multiplier m53(A[address][21],B[21][1],mul53);   multiplier m54(A[address][22],B[22][1],mul54);   multiplier m55(A[address][23],B[23][1],mul55);   multiplier m56(A[address][24],B[24][1],mul56);   multiplier m57(A[address][25],B[25][1],mul57);   multiplier m58(A[address][26],B[26][1],mul58);   multiplier m59(A[address][27],B[27][1],mul59);   multiplier m60(A[address][28],B[28][1],mul60);   multiplier m61(A[address][29],B[29][1],mul61);   multiplier m62(A[address][30],B[30][1],mul62);   multiplier m63(A[address][31],B[31][1],mul63);   
	multiplier m64(A[address][0],B[0][2],mul64);   multiplier m65(A[address][1],B[1][2],mul65);   multiplier m66(A[address][2],B[2][2],mul66);   multiplier m67(A[address][3],B[3][2],mul67);   multiplier m68(A[address][4],B[4][2],mul68);   multiplier m69(A[address][5],B[5][2],mul69);   multiplier m70(A[address][6],B[6][2],mul70);   multiplier m71(A[address][7],B[7][2],mul71);   multiplier m72(A[address][8],B[8][2],mul72);   multiplier m73(A[address][9],B[9][2],mul73);   multiplier m74(A[address][10],B[10][2],mul74);   multiplier m75(A[address][11],B[11][2],mul75);   multiplier m76(A[address][12],B[12][2],mul76);   multiplier m77(A[address][13],B[13][2],mul77);   multiplier m78(A[address][14],B[14][2],mul78);   multiplier m79(A[address][15],B[15][2],mul79);   multiplier m80(A[address][16],B[16][2],mul80);   multiplier m81(A[address][17],B[17][2],mul81);   multiplier m82(A[address][18],B[18][2],mul82);   multiplier m83(A[address][19],B[19][2],mul83);   multiplier m84(A[address][20],B[20][2],mul84);   multiplier m85(A[address][21],B[21][2],mul85);   multiplier m86(A[address][22],B[22][2],mul86);   multiplier m87(A[address][23],B[23][2],mul87);   multiplier m88(A[address][24],B[24][2],mul88);   multiplier m89(A[address][25],B[25][2],mul89);   multiplier m90(A[address][26],B[26][2],mul90);   multiplier m91(A[address][27],B[27][2],mul91);   multiplier m92(A[address][28],B[28][2],mul92);   multiplier m93(A[address][29],B[29][2],mul93);   multiplier m94(A[address][30],B[30][2],mul94);   multiplier m95(A[address][31],B[31][2],mul95);   
	multiplier m96(A[address][0],B[0][3],mul96);   multiplier m97(A[address][1],B[1][3],mul97);   multiplier m98(A[address][2],B[2][3],mul98);   multiplier m99(A[address][3],B[3][3],mul99);   multiplier m100(A[address][4],B[4][3],mul100);   multiplier m101(A[address][5],B[5][3],mul101);   multiplier m102(A[address][6],B[6][3],mul102);   multiplier m103(A[address][7],B[7][3],mul103);   multiplier m104(A[address][8],B[8][3],mul104);   multiplier m105(A[address][9],B[9][3],mul105);   multiplier m106(A[address][10],B[10][3],mul106);   multiplier m107(A[address][11],B[11][3],mul107);   multiplier m108(A[address][12],B[12][3],mul108);   multiplier m109(A[address][13],B[13][3],mul109);   multiplier m110(A[address][14],B[14][3],mul110);   multiplier m111(A[address][15],B[15][3],mul111);   multiplier m112(A[address][16],B[16][3],mul112);   multiplier m113(A[address][17],B[17][3],mul113);   multiplier m114(A[address][18],B[18][3],mul114);   multiplier m115(A[address][19],B[19][3],mul115);   multiplier m116(A[address][20],B[20][3],mul116);   multiplier m117(A[address][21],B[21][3],mul117);   multiplier m118(A[address][22],B[22][3],mul118);   multiplier m119(A[address][23],B[23][3],mul119);   multiplier m120(A[address][24],B[24][3],mul120);   multiplier m121(A[address][25],B[25][3],mul121);   multiplier m122(A[address][26],B[26][3],mul122);   multiplier m123(A[address][27],B[27][3],mul123);   multiplier m124(A[address][28],B[28][3],mul124);   multiplier m125(A[address][29],B[29][3],mul125);   multiplier m126(A[address][30],B[30][3],mul126);   multiplier m127(A[address][31],B[31][3],mul127);   
	multiplier m128(A[address][0],B[0][4],mul128);   multiplier m129(A[address][1],B[1][4],mul129);   multiplier m130(A[address][2],B[2][4],mul130);   multiplier m131(A[address][3],B[3][4],mul131);   multiplier m132(A[address][4],B[4][4],mul132);   multiplier m133(A[address][5],B[5][4],mul133);   multiplier m134(A[address][6],B[6][4],mul134);   multiplier m135(A[address][7],B[7][4],mul135);   multiplier m136(A[address][8],B[8][4],mul136);   multiplier m137(A[address][9],B[9][4],mul137);   multiplier m138(A[address][10],B[10][4],mul138);   multiplier m139(A[address][11],B[11][4],mul139);   multiplier m140(A[address][12],B[12][4],mul140);   multiplier m141(A[address][13],B[13][4],mul141);   multiplier m142(A[address][14],B[14][4],mul142);   multiplier m143(A[address][15],B[15][4],mul143);   multiplier m144(A[address][16],B[16][4],mul144);   multiplier m145(A[address][17],B[17][4],mul145);   multiplier m146(A[address][18],B[18][4],mul146);   multiplier m147(A[address][19],B[19][4],mul147);   multiplier m148(A[address][20],B[20][4],mul148);   multiplier m149(A[address][21],B[21][4],mul149);   multiplier m150(A[address][22],B[22][4],mul150);   multiplier m151(A[address][23],B[23][4],mul151);   multiplier m152(A[address][24],B[24][4],mul152);   multiplier m153(A[address][25],B[25][4],mul153);   multiplier m154(A[address][26],B[26][4],mul154);   multiplier m155(A[address][27],B[27][4],mul155);   multiplier m156(A[address][28],B[28][4],mul156);   multiplier m157(A[address][29],B[29][4],mul157);   multiplier m158(A[address][30],B[30][4],mul158);   multiplier m159(A[address][31],B[31][4],mul159);   
	multiplier m160(A[address][0],B[0][5],mul160);   multiplier m161(A[address][1],B[1][5],mul161);   multiplier m162(A[address][2],B[2][5],mul162);   multiplier m163(A[address][3],B[3][5],mul163);   multiplier m164(A[address][4],B[4][5],mul164);   multiplier m165(A[address][5],B[5][5],mul165);   multiplier m166(A[address][6],B[6][5],mul166);   multiplier m167(A[address][7],B[7][5],mul167);   multiplier m168(A[address][8],B[8][5],mul168);   multiplier m169(A[address][9],B[9][5],mul169);   multiplier m170(A[address][10],B[10][5],mul170);   multiplier m171(A[address][11],B[11][5],mul171);   multiplier m172(A[address][12],B[12][5],mul172);   multiplier m173(A[address][13],B[13][5],mul173);   multiplier m174(A[address][14],B[14][5],mul174);   multiplier m175(A[address][15],B[15][5],mul175);   multiplier m176(A[address][16],B[16][5],mul176);   multiplier m177(A[address][17],B[17][5],mul177);   multiplier m178(A[address][18],B[18][5],mul178);   multiplier m179(A[address][19],B[19][5],mul179);   multiplier m180(A[address][20],B[20][5],mul180);   multiplier m181(A[address][21],B[21][5],mul181);   multiplier m182(A[address][22],B[22][5],mul182);   multiplier m183(A[address][23],B[23][5],mul183);   multiplier m184(A[address][24],B[24][5],mul184);   multiplier m185(A[address][25],B[25][5],mul185);   multiplier m186(A[address][26],B[26][5],mul186);   multiplier m187(A[address][27],B[27][5],mul187);   multiplier m188(A[address][28],B[28][5],mul188);   multiplier m189(A[address][29],B[29][5],mul189);   multiplier m190(A[address][30],B[30][5],mul190);   multiplier m191(A[address][31],B[31][5],mul191);   
	multiplier m192(A[address][0],B[0][6],mul192);   multiplier m193(A[address][1],B[1][6],mul193);   multiplier m194(A[address][2],B[2][6],mul194);   multiplier m195(A[address][3],B[3][6],mul195);   multiplier m196(A[address][4],B[4][6],mul196);   multiplier m197(A[address][5],B[5][6],mul197);   multiplier m198(A[address][6],B[6][6],mul198);   multiplier m199(A[address][7],B[7][6],mul199);   multiplier m200(A[address][8],B[8][6],mul200);   multiplier m201(A[address][9],B[9][6],mul201);   multiplier m202(A[address][10],B[10][6],mul202);   multiplier m203(A[address][11],B[11][6],mul203);   multiplier m204(A[address][12],B[12][6],mul204);   multiplier m205(A[address][13],B[13][6],mul205);   multiplier m206(A[address][14],B[14][6],mul206);   multiplier m207(A[address][15],B[15][6],mul207);   multiplier m208(A[address][16],B[16][6],mul208);   multiplier m209(A[address][17],B[17][6],mul209);   multiplier m210(A[address][18],B[18][6],mul210);   multiplier m211(A[address][19],B[19][6],mul211);   multiplier m212(A[address][20],B[20][6],mul212);   multiplier m213(A[address][21],B[21][6],mul213);   multiplier m214(A[address][22],B[22][6],mul214);   multiplier m215(A[address][23],B[23][6],mul215);   multiplier m216(A[address][24],B[24][6],mul216);   multiplier m217(A[address][25],B[25][6],mul217);   multiplier m218(A[address][26],B[26][6],mul218);   multiplier m219(A[address][27],B[27][6],mul219);   multiplier m220(A[address][28],B[28][6],mul220);   multiplier m221(A[address][29],B[29][6],mul221);   multiplier m222(A[address][30],B[30][6],mul222);   multiplier m223(A[address][31],B[31][6],mul223);   
	multiplier m224(A[address][0],B[0][7],mul224);   multiplier m225(A[address][1],B[1][7],mul225);   multiplier m226(A[address][2],B[2][7],mul226);   multiplier m227(A[address][3],B[3][7],mul227);   multiplier m228(A[address][4],B[4][7],mul228);   multiplier m229(A[address][5],B[5][7],mul229);   multiplier m230(A[address][6],B[6][7],mul230);   multiplier m231(A[address][7],B[7][7],mul231);   multiplier m232(A[address][8],B[8][7],mul232);   multiplier m233(A[address][9],B[9][7],mul233);   multiplier m234(A[address][10],B[10][7],mul234);   multiplier m235(A[address][11],B[11][7],mul235);   multiplier m236(A[address][12],B[12][7],mul236);   multiplier m237(A[address][13],B[13][7],mul237);   multiplier m238(A[address][14],B[14][7],mul238);   multiplier m239(A[address][15],B[15][7],mul239);   multiplier m240(A[address][16],B[16][7],mul240);   multiplier m241(A[address][17],B[17][7],mul241);   multiplier m242(A[address][18],B[18][7],mul242);   multiplier m243(A[address][19],B[19][7],mul243);   multiplier m244(A[address][20],B[20][7],mul244);   multiplier m245(A[address][21],B[21][7],mul245);   multiplier m246(A[address][22],B[22][7],mul246);   multiplier m247(A[address][23],B[23][7],mul247);   multiplier m248(A[address][24],B[24][7],mul248);   multiplier m249(A[address][25],B[25][7],mul249);   multiplier m250(A[address][26],B[26][7],mul250);   multiplier m251(A[address][27],B[27][7],mul251);   multiplier m252(A[address][28],B[28][7],mul252);   multiplier m253(A[address][29],B[29][7],mul253);   multiplier m254(A[address][30],B[30][7],mul254);   multiplier m255(A[address][31],B[31][7],mul255);   
	multiplier m256(A[address][0],B[0][8],mul256);   multiplier m257(A[address][1],B[1][8],mul257);   multiplier m258(A[address][2],B[2][8],mul258);   multiplier m259(A[address][3],B[3][8],mul259);   multiplier m260(A[address][4],B[4][8],mul260);   multiplier m261(A[address][5],B[5][8],mul261);   multiplier m262(A[address][6],B[6][8],mul262);   multiplier m263(A[address][7],B[7][8],mul263);   multiplier m264(A[address][8],B[8][8],mul264);   multiplier m265(A[address][9],B[9][8],mul265);   multiplier m266(A[address][10],B[10][8],mul266);   multiplier m267(A[address][11],B[11][8],mul267);   multiplier m268(A[address][12],B[12][8],mul268);   multiplier m269(A[address][13],B[13][8],mul269);   multiplier m270(A[address][14],B[14][8],mul270);   multiplier m271(A[address][15],B[15][8],mul271);   multiplier m272(A[address][16],B[16][8],mul272);   multiplier m273(A[address][17],B[17][8],mul273);   multiplier m274(A[address][18],B[18][8],mul274);   multiplier m275(A[address][19],B[19][8],mul275);   multiplier m276(A[address][20],B[20][8],mul276);   multiplier m277(A[address][21],B[21][8],mul277);   multiplier m278(A[address][22],B[22][8],mul278);   multiplier m279(A[address][23],B[23][8],mul279);   multiplier m280(A[address][24],B[24][8],mul280);   multiplier m281(A[address][25],B[25][8],mul281);   multiplier m282(A[address][26],B[26][8],mul282);   multiplier m283(A[address][27],B[27][8],mul283);   multiplier m284(A[address][28],B[28][8],mul284);   multiplier m285(A[address][29],B[29][8],mul285);   multiplier m286(A[address][30],B[30][8],mul286);   multiplier m287(A[address][31],B[31][8],mul287);   
	multiplier m288(A[address][0],B[0][9],mul288);   multiplier m289(A[address][1],B[1][9],mul289);   multiplier m290(A[address][2],B[2][9],mul290);   multiplier m291(A[address][3],B[3][9],mul291);   multiplier m292(A[address][4],B[4][9],mul292);   multiplier m293(A[address][5],B[5][9],mul293);   multiplier m294(A[address][6],B[6][9],mul294);   multiplier m295(A[address][7],B[7][9],mul295);   multiplier m296(A[address][8],B[8][9],mul296);   multiplier m297(A[address][9],B[9][9],mul297);   multiplier m298(A[address][10],B[10][9],mul298);   multiplier m299(A[address][11],B[11][9],mul299);   multiplier m300(A[address][12],B[12][9],mul300);   multiplier m301(A[address][13],B[13][9],mul301);   multiplier m302(A[address][14],B[14][9],mul302);   multiplier m303(A[address][15],B[15][9],mul303);   multiplier m304(A[address][16],B[16][9],mul304);   multiplier m305(A[address][17],B[17][9],mul305);   multiplier m306(A[address][18],B[18][9],mul306);   multiplier m307(A[address][19],B[19][9],mul307);   multiplier m308(A[address][20],B[20][9],mul308);   multiplier m309(A[address][21],B[21][9],mul309);   multiplier m310(A[address][22],B[22][9],mul310);   multiplier m311(A[address][23],B[23][9],mul311);   multiplier m312(A[address][24],B[24][9],mul312);   multiplier m313(A[address][25],B[25][9],mul313);   multiplier m314(A[address][26],B[26][9],mul314);   multiplier m315(A[address][27],B[27][9],mul315);   multiplier m316(A[address][28],B[28][9],mul316);   multiplier m317(A[address][29],B[29][9],mul317);   multiplier m318(A[address][30],B[30][9],mul318);   multiplier m319(A[address][31],B[31][9],mul319);   
	multiplier m320(A[address][0],B[0][10],mul320);   multiplier m321(A[address][1],B[1][10],mul321);   multiplier m322(A[address][2],B[2][10],mul322);   multiplier m323(A[address][3],B[3][10],mul323);   multiplier m324(A[address][4],B[4][10],mul324);   multiplier m325(A[address][5],B[5][10],mul325);   multiplier m326(A[address][6],B[6][10],mul326);   multiplier m327(A[address][7],B[7][10],mul327);   multiplier m328(A[address][8],B[8][10],mul328);   multiplier m329(A[address][9],B[9][10],mul329);   multiplier m330(A[address][10],B[10][10],mul330);   multiplier m331(A[address][11],B[11][10],mul331);   multiplier m332(A[address][12],B[12][10],mul332);   multiplier m333(A[address][13],B[13][10],mul333);   multiplier m334(A[address][14],B[14][10],mul334);   multiplier m335(A[address][15],B[15][10],mul335);   multiplier m336(A[address][16],B[16][10],mul336);   multiplier m337(A[address][17],B[17][10],mul337);   multiplier m338(A[address][18],B[18][10],mul338);   multiplier m339(A[address][19],B[19][10],mul339);   multiplier m340(A[address][20],B[20][10],mul340);   multiplier m341(A[address][21],B[21][10],mul341);   multiplier m342(A[address][22],B[22][10],mul342);   multiplier m343(A[address][23],B[23][10],mul343);   multiplier m344(A[address][24],B[24][10],mul344);   multiplier m345(A[address][25],B[25][10],mul345);   multiplier m346(A[address][26],B[26][10],mul346);   multiplier m347(A[address][27],B[27][10],mul347);   multiplier m348(A[address][28],B[28][10],mul348);   multiplier m349(A[address][29],B[29][10],mul349);   multiplier m350(A[address][30],B[30][10],mul350);   multiplier m351(A[address][31],B[31][10],mul351);   
	multiplier m352(A[address][0],B[0][11],mul352);   multiplier m353(A[address][1],B[1][11],mul353);   multiplier m354(A[address][2],B[2][11],mul354);   multiplier m355(A[address][3],B[3][11],mul355);   multiplier m356(A[address][4],B[4][11],mul356);   multiplier m357(A[address][5],B[5][11],mul357);   multiplier m358(A[address][6],B[6][11],mul358);   multiplier m359(A[address][7],B[7][11],mul359);   multiplier m360(A[address][8],B[8][11],mul360);   multiplier m361(A[address][9],B[9][11],mul361);   multiplier m362(A[address][10],B[10][11],mul362);   multiplier m363(A[address][11],B[11][11],mul363);   multiplier m364(A[address][12],B[12][11],mul364);   multiplier m365(A[address][13],B[13][11],mul365);   multiplier m366(A[address][14],B[14][11],mul366);   multiplier m367(A[address][15],B[15][11],mul367);   multiplier m368(A[address][16],B[16][11],mul368);   multiplier m369(A[address][17],B[17][11],mul369);   multiplier m370(A[address][18],B[18][11],mul370);   multiplier m371(A[address][19],B[19][11],mul371);   multiplier m372(A[address][20],B[20][11],mul372);   multiplier m373(A[address][21],B[21][11],mul373);   multiplier m374(A[address][22],B[22][11],mul374);   multiplier m375(A[address][23],B[23][11],mul375);   multiplier m376(A[address][24],B[24][11],mul376);   multiplier m377(A[address][25],B[25][11],mul377);   multiplier m378(A[address][26],B[26][11],mul378);   multiplier m379(A[address][27],B[27][11],mul379);   multiplier m380(A[address][28],B[28][11],mul380);   multiplier m381(A[address][29],B[29][11],mul381);   multiplier m382(A[address][30],B[30][11],mul382);   multiplier m383(A[address][31],B[31][11],mul383);   
	multiplier m384(A[address][0],B[0][12],mul384);   multiplier m385(A[address][1],B[1][12],mul385);   multiplier m386(A[address][2],B[2][12],mul386);   multiplier m387(A[address][3],B[3][12],mul387);   multiplier m388(A[address][4],B[4][12],mul388);   multiplier m389(A[address][5],B[5][12],mul389);   multiplier m390(A[address][6],B[6][12],mul390);   multiplier m391(A[address][7],B[7][12],mul391);   multiplier m392(A[address][8],B[8][12],mul392);   multiplier m393(A[address][9],B[9][12],mul393);   multiplier m394(A[address][10],B[10][12],mul394);   multiplier m395(A[address][11],B[11][12],mul395);   multiplier m396(A[address][12],B[12][12],mul396);   multiplier m397(A[address][13],B[13][12],mul397);   multiplier m398(A[address][14],B[14][12],mul398);   multiplier m399(A[address][15],B[15][12],mul399);   multiplier m400(A[address][16],B[16][12],mul400);   multiplier m401(A[address][17],B[17][12],mul401);   multiplier m402(A[address][18],B[18][12],mul402);   multiplier m403(A[address][19],B[19][12],mul403);   multiplier m404(A[address][20],B[20][12],mul404);   multiplier m405(A[address][21],B[21][12],mul405);   multiplier m406(A[address][22],B[22][12],mul406);   multiplier m407(A[address][23],B[23][12],mul407);   multiplier m408(A[address][24],B[24][12],mul408);   multiplier m409(A[address][25],B[25][12],mul409);   multiplier m410(A[address][26],B[26][12],mul410);   multiplier m411(A[address][27],B[27][12],mul411);   multiplier m412(A[address][28],B[28][12],mul412);   multiplier m413(A[address][29],B[29][12],mul413);   multiplier m414(A[address][30],B[30][12],mul414);   multiplier m415(A[address][31],B[31][12],mul415);   
	multiplier m416(A[address][0],B[0][13],mul416);   multiplier m417(A[address][1],B[1][13],mul417);   multiplier m418(A[address][2],B[2][13],mul418);   multiplier m419(A[address][3],B[3][13],mul419);   multiplier m420(A[address][4],B[4][13],mul420);   multiplier m421(A[address][5],B[5][13],mul421);   multiplier m422(A[address][6],B[6][13],mul422);   multiplier m423(A[address][7],B[7][13],mul423);   multiplier m424(A[address][8],B[8][13],mul424);   multiplier m425(A[address][9],B[9][13],mul425);   multiplier m426(A[address][10],B[10][13],mul426);   multiplier m427(A[address][11],B[11][13],mul427);   multiplier m428(A[address][12],B[12][13],mul428);   multiplier m429(A[address][13],B[13][13],mul429);   multiplier m430(A[address][14],B[14][13],mul430);   multiplier m431(A[address][15],B[15][13],mul431);   multiplier m432(A[address][16],B[16][13],mul432);   multiplier m433(A[address][17],B[17][13],mul433);   multiplier m434(A[address][18],B[18][13],mul434);   multiplier m435(A[address][19],B[19][13],mul435);   multiplier m436(A[address][20],B[20][13],mul436);   multiplier m437(A[address][21],B[21][13],mul437);   multiplier m438(A[address][22],B[22][13],mul438);   multiplier m439(A[address][23],B[23][13],mul439);   multiplier m440(A[address][24],B[24][13],mul440);   multiplier m441(A[address][25],B[25][13],mul441);   multiplier m442(A[address][26],B[26][13],mul442);   multiplier m443(A[address][27],B[27][13],mul443);   multiplier m444(A[address][28],B[28][13],mul444);   multiplier m445(A[address][29],B[29][13],mul445);   multiplier m446(A[address][30],B[30][13],mul446);   multiplier m447(A[address][31],B[31][13],mul447);   
	multiplier m448(A[address][0],B[0][14],mul448);   multiplier m449(A[address][1],B[1][14],mul449);   multiplier m450(A[address][2],B[2][14],mul450);   multiplier m451(A[address][3],B[3][14],mul451);   multiplier m452(A[address][4],B[4][14],mul452);   multiplier m453(A[address][5],B[5][14],mul453);   multiplier m454(A[address][6],B[6][14],mul454);   multiplier m455(A[address][7],B[7][14],mul455);   multiplier m456(A[address][8],B[8][14],mul456);   multiplier m457(A[address][9],B[9][14],mul457);   multiplier m458(A[address][10],B[10][14],mul458);   multiplier m459(A[address][11],B[11][14],mul459);   multiplier m460(A[address][12],B[12][14],mul460);   multiplier m461(A[address][13],B[13][14],mul461);   multiplier m462(A[address][14],B[14][14],mul462);   multiplier m463(A[address][15],B[15][14],mul463);   multiplier m464(A[address][16],B[16][14],mul464);   multiplier m465(A[address][17],B[17][14],mul465);   multiplier m466(A[address][18],B[18][14],mul466);   multiplier m467(A[address][19],B[19][14],mul467);   multiplier m468(A[address][20],B[20][14],mul468);   multiplier m469(A[address][21],B[21][14],mul469);   multiplier m470(A[address][22],B[22][14],mul470);   multiplier m471(A[address][23],B[23][14],mul471);   multiplier m472(A[address][24],B[24][14],mul472);   multiplier m473(A[address][25],B[25][14],mul473);   multiplier m474(A[address][26],B[26][14],mul474);   multiplier m475(A[address][27],B[27][14],mul475);   multiplier m476(A[address][28],B[28][14],mul476);   multiplier m477(A[address][29],B[29][14],mul477);   multiplier m478(A[address][30],B[30][14],mul478);   multiplier m479(A[address][31],B[31][14],mul479);   
	multiplier m480(A[address][0],B[0][15],mul480);   multiplier m481(A[address][1],B[1][15],mul481);   multiplier m482(A[address][2],B[2][15],mul482);   multiplier m483(A[address][3],B[3][15],mul483);   multiplier m484(A[address][4],B[4][15],mul484);   multiplier m485(A[address][5],B[5][15],mul485);   multiplier m486(A[address][6],B[6][15],mul486);   multiplier m487(A[address][7],B[7][15],mul487);   multiplier m488(A[address][8],B[8][15],mul488);   multiplier m489(A[address][9],B[9][15],mul489);   multiplier m490(A[address][10],B[10][15],mul490);   multiplier m491(A[address][11],B[11][15],mul491);   multiplier m492(A[address][12],B[12][15],mul492);   multiplier m493(A[address][13],B[13][15],mul493);   multiplier m494(A[address][14],B[14][15],mul494);   multiplier m495(A[address][15],B[15][15],mul495);   multiplier m496(A[address][16],B[16][15],mul496);   multiplier m497(A[address][17],B[17][15],mul497);   multiplier m498(A[address][18],B[18][15],mul498);   multiplier m499(A[address][19],B[19][15],mul499);   multiplier m500(A[address][20],B[20][15],mul500);   multiplier m501(A[address][21],B[21][15],mul501);   multiplier m502(A[address][22],B[22][15],mul502);   multiplier m503(A[address][23],B[23][15],mul503);   multiplier m504(A[address][24],B[24][15],mul504);   multiplier m505(A[address][25],B[25][15],mul505);   multiplier m506(A[address][26],B[26][15],mul506);   multiplier m507(A[address][27],B[27][15],mul507);   multiplier m508(A[address][28],B[28][15],mul508);   multiplier m509(A[address][29],B[29][15],mul509);   multiplier m510(A[address][30],B[30][15],mul510);   multiplier m511(A[address][31],B[31][15],mul511);   
	multiplier m512(A[address][0],B[0][16],mul512);   multiplier m513(A[address][1],B[1][16],mul513);   multiplier m514(A[address][2],B[2][16],mul514);   multiplier m515(A[address][3],B[3][16],mul515);   multiplier m516(A[address][4],B[4][16],mul516);   multiplier m517(A[address][5],B[5][16],mul517);   multiplier m518(A[address][6],B[6][16],mul518);   multiplier m519(A[address][7],B[7][16],mul519);   multiplier m520(A[address][8],B[8][16],mul520);   multiplier m521(A[address][9],B[9][16],mul521);   multiplier m522(A[address][10],B[10][16],mul522);   multiplier m523(A[address][11],B[11][16],mul523);   multiplier m524(A[address][12],B[12][16],mul524);   multiplier m525(A[address][13],B[13][16],mul525);   multiplier m526(A[address][14],B[14][16],mul526);   multiplier m527(A[address][15],B[15][16],mul527);   multiplier m528(A[address][16],B[16][16],mul528);   multiplier m529(A[address][17],B[17][16],mul529);   multiplier m530(A[address][18],B[18][16],mul530);   multiplier m531(A[address][19],B[19][16],mul531);   multiplier m532(A[address][20],B[20][16],mul532);   multiplier m533(A[address][21],B[21][16],mul533);   multiplier m534(A[address][22],B[22][16],mul534);   multiplier m535(A[address][23],B[23][16],mul535);   multiplier m536(A[address][24],B[24][16],mul536);   multiplier m537(A[address][25],B[25][16],mul537);   multiplier m538(A[address][26],B[26][16],mul538);   multiplier m539(A[address][27],B[27][16],mul539);   multiplier m540(A[address][28],B[28][16],mul540);   multiplier m541(A[address][29],B[29][16],mul541);   multiplier m542(A[address][30],B[30][16],mul542);   multiplier m543(A[address][31],B[31][16],mul543);   
	multiplier m544(A[address][0],B[0][17],mul544);   multiplier m545(A[address][1],B[1][17],mul545);   multiplier m546(A[address][2],B[2][17],mul546);   multiplier m547(A[address][3],B[3][17],mul547);   multiplier m548(A[address][4],B[4][17],mul548);   multiplier m549(A[address][5],B[5][17],mul549);   multiplier m550(A[address][6],B[6][17],mul550);   multiplier m551(A[address][7],B[7][17],mul551);   multiplier m552(A[address][8],B[8][17],mul552);   multiplier m553(A[address][9],B[9][17],mul553);   multiplier m554(A[address][10],B[10][17],mul554);   multiplier m555(A[address][11],B[11][17],mul555);   multiplier m556(A[address][12],B[12][17],mul556);   multiplier m557(A[address][13],B[13][17],mul557);   multiplier m558(A[address][14],B[14][17],mul558);   multiplier m559(A[address][15],B[15][17],mul559);   multiplier m560(A[address][16],B[16][17],mul560);   multiplier m561(A[address][17],B[17][17],mul561);   multiplier m562(A[address][18],B[18][17],mul562);   multiplier m563(A[address][19],B[19][17],mul563);   multiplier m564(A[address][20],B[20][17],mul564);   multiplier m565(A[address][21],B[21][17],mul565);   multiplier m566(A[address][22],B[22][17],mul566);   multiplier m567(A[address][23],B[23][17],mul567);   multiplier m568(A[address][24],B[24][17],mul568);   multiplier m569(A[address][25],B[25][17],mul569);   multiplier m570(A[address][26],B[26][17],mul570);   multiplier m571(A[address][27],B[27][17],mul571);   multiplier m572(A[address][28],B[28][17],mul572);   multiplier m573(A[address][29],B[29][17],mul573);   multiplier m574(A[address][30],B[30][17],mul574);   multiplier m575(A[address][31],B[31][17],mul575);   
	multiplier m576(A[address][0],B[0][18],mul576);   multiplier m577(A[address][1],B[1][18],mul577);   multiplier m578(A[address][2],B[2][18],mul578);   multiplier m579(A[address][3],B[3][18],mul579);   multiplier m580(A[address][4],B[4][18],mul580);   multiplier m581(A[address][5],B[5][18],mul581);   multiplier m582(A[address][6],B[6][18],mul582);   multiplier m583(A[address][7],B[7][18],mul583);   multiplier m584(A[address][8],B[8][18],mul584);   multiplier m585(A[address][9],B[9][18],mul585);   multiplier m586(A[address][10],B[10][18],mul586);   multiplier m587(A[address][11],B[11][18],mul587);   multiplier m588(A[address][12],B[12][18],mul588);   multiplier m589(A[address][13],B[13][18],mul589);   multiplier m590(A[address][14],B[14][18],mul590);   multiplier m591(A[address][15],B[15][18],mul591);   multiplier m592(A[address][16],B[16][18],mul592);   multiplier m593(A[address][17],B[17][18],mul593);   multiplier m594(A[address][18],B[18][18],mul594);   multiplier m595(A[address][19],B[19][18],mul595);   multiplier m596(A[address][20],B[20][18],mul596);   multiplier m597(A[address][21],B[21][18],mul597);   multiplier m598(A[address][22],B[22][18],mul598);   multiplier m599(A[address][23],B[23][18],mul599);   multiplier m600(A[address][24],B[24][18],mul600);   multiplier m601(A[address][25],B[25][18],mul601);   multiplier m602(A[address][26],B[26][18],mul602);   multiplier m603(A[address][27],B[27][18],mul603);   multiplier m604(A[address][28],B[28][18],mul604);   multiplier m605(A[address][29],B[29][18],mul605);   multiplier m606(A[address][30],B[30][18],mul606);   multiplier m607(A[address][31],B[31][18],mul607);   
	multiplier m608(A[address][0],B[0][19],mul608);   multiplier m609(A[address][1],B[1][19],mul609);   multiplier m610(A[address][2],B[2][19],mul610);   multiplier m611(A[address][3],B[3][19],mul611);   multiplier m612(A[address][4],B[4][19],mul612);   multiplier m613(A[address][5],B[5][19],mul613);   multiplier m614(A[address][6],B[6][19],mul614);   multiplier m615(A[address][7],B[7][19],mul615);   multiplier m616(A[address][8],B[8][19],mul616);   multiplier m617(A[address][9],B[9][19],mul617);   multiplier m618(A[address][10],B[10][19],mul618);   multiplier m619(A[address][11],B[11][19],mul619);   multiplier m620(A[address][12],B[12][19],mul620);   multiplier m621(A[address][13],B[13][19],mul621);   multiplier m622(A[address][14],B[14][19],mul622);   multiplier m623(A[address][15],B[15][19],mul623);   multiplier m624(A[address][16],B[16][19],mul624);   multiplier m625(A[address][17],B[17][19],mul625);   multiplier m626(A[address][18],B[18][19],mul626);   multiplier m627(A[address][19],B[19][19],mul627);   multiplier m628(A[address][20],B[20][19],mul628);   multiplier m629(A[address][21],B[21][19],mul629);   multiplier m630(A[address][22],B[22][19],mul630);   multiplier m631(A[address][23],B[23][19],mul631);   multiplier m632(A[address][24],B[24][19],mul632);   multiplier m633(A[address][25],B[25][19],mul633);   multiplier m634(A[address][26],B[26][19],mul634);   multiplier m635(A[address][27],B[27][19],mul635);   multiplier m636(A[address][28],B[28][19],mul636);   multiplier m637(A[address][29],B[29][19],mul637);   multiplier m638(A[address][30],B[30][19],mul638);   multiplier m639(A[address][31],B[31][19],mul639);   
	multiplier m640(A[address][0],B[0][20],mul640);   multiplier m641(A[address][1],B[1][20],mul641);   multiplier m642(A[address][2],B[2][20],mul642);   multiplier m643(A[address][3],B[3][20],mul643);   multiplier m644(A[address][4],B[4][20],mul644);   multiplier m645(A[address][5],B[5][20],mul645);   multiplier m646(A[address][6],B[6][20],mul646);   multiplier m647(A[address][7],B[7][20],mul647);   multiplier m648(A[address][8],B[8][20],mul648);   multiplier m649(A[address][9],B[9][20],mul649);   multiplier m650(A[address][10],B[10][20],mul650);   multiplier m651(A[address][11],B[11][20],mul651);   multiplier m652(A[address][12],B[12][20],mul652);   multiplier m653(A[address][13],B[13][20],mul653);   multiplier m654(A[address][14],B[14][20],mul654);   multiplier m655(A[address][15],B[15][20],mul655);   multiplier m656(A[address][16],B[16][20],mul656);   multiplier m657(A[address][17],B[17][20],mul657);   multiplier m658(A[address][18],B[18][20],mul658);   multiplier m659(A[address][19],B[19][20],mul659);   multiplier m660(A[address][20],B[20][20],mul660);   multiplier m661(A[address][21],B[21][20],mul661);   multiplier m662(A[address][22],B[22][20],mul662);   multiplier m663(A[address][23],B[23][20],mul663);   multiplier m664(A[address][24],B[24][20],mul664);   multiplier m665(A[address][25],B[25][20],mul665);   multiplier m666(A[address][26],B[26][20],mul666);   multiplier m667(A[address][27],B[27][20],mul667);   multiplier m668(A[address][28],B[28][20],mul668);   multiplier m669(A[address][29],B[29][20],mul669);   multiplier m670(A[address][30],B[30][20],mul670);   multiplier m671(A[address][31],B[31][20],mul671);   
	multiplier m672(A[address][0],B[0][21],mul672);   multiplier m673(A[address][1],B[1][21],mul673);   multiplier m674(A[address][2],B[2][21],mul674);   multiplier m675(A[address][3],B[3][21],mul675);   multiplier m676(A[address][4],B[4][21],mul676);   multiplier m677(A[address][5],B[5][21],mul677);   multiplier m678(A[address][6],B[6][21],mul678);   multiplier m679(A[address][7],B[7][21],mul679);   multiplier m680(A[address][8],B[8][21],mul680);   multiplier m681(A[address][9],B[9][21],mul681);   multiplier m682(A[address][10],B[10][21],mul682);   multiplier m683(A[address][11],B[11][21],mul683);   multiplier m684(A[address][12],B[12][21],mul684);   multiplier m685(A[address][13],B[13][21],mul685);   multiplier m686(A[address][14],B[14][21],mul686);   multiplier m687(A[address][15],B[15][21],mul687);   multiplier m688(A[address][16],B[16][21],mul688);   multiplier m689(A[address][17],B[17][21],mul689);   multiplier m690(A[address][18],B[18][21],mul690);   multiplier m691(A[address][19],B[19][21],mul691);   multiplier m692(A[address][20],B[20][21],mul692);   multiplier m693(A[address][21],B[21][21],mul693);   multiplier m694(A[address][22],B[22][21],mul694);   multiplier m695(A[address][23],B[23][21],mul695);   multiplier m696(A[address][24],B[24][21],mul696);   multiplier m697(A[address][25],B[25][21],mul697);   multiplier m698(A[address][26],B[26][21],mul698);   multiplier m699(A[address][27],B[27][21],mul699);   multiplier m700(A[address][28],B[28][21],mul700);   multiplier m701(A[address][29],B[29][21],mul701);   multiplier m702(A[address][30],B[30][21],mul702);   multiplier m703(A[address][31],B[31][21],mul703);   
	multiplier m704(A[address][0],B[0][22],mul704);   multiplier m705(A[address][1],B[1][22],mul705);   multiplier m706(A[address][2],B[2][22],mul706);   multiplier m707(A[address][3],B[3][22],mul707);   multiplier m708(A[address][4],B[4][22],mul708);   multiplier m709(A[address][5],B[5][22],mul709);   multiplier m710(A[address][6],B[6][22],mul710);   multiplier m711(A[address][7],B[7][22],mul711);   multiplier m712(A[address][8],B[8][22],mul712);   multiplier m713(A[address][9],B[9][22],mul713);   multiplier m714(A[address][10],B[10][22],mul714);   multiplier m715(A[address][11],B[11][22],mul715);   multiplier m716(A[address][12],B[12][22],mul716);   multiplier m717(A[address][13],B[13][22],mul717);   multiplier m718(A[address][14],B[14][22],mul718);   multiplier m719(A[address][15],B[15][22],mul719);   multiplier m720(A[address][16],B[16][22],mul720);   multiplier m721(A[address][17],B[17][22],mul721);   multiplier m722(A[address][18],B[18][22],mul722);   multiplier m723(A[address][19],B[19][22],mul723);   multiplier m724(A[address][20],B[20][22],mul724);   multiplier m725(A[address][21],B[21][22],mul725);   multiplier m726(A[address][22],B[22][22],mul726);   multiplier m727(A[address][23],B[23][22],mul727);   multiplier m728(A[address][24],B[24][22],mul728);   multiplier m729(A[address][25],B[25][22],mul729);   multiplier m730(A[address][26],B[26][22],mul730);   multiplier m731(A[address][27],B[27][22],mul731);   multiplier m732(A[address][28],B[28][22],mul732);   multiplier m733(A[address][29],B[29][22],mul733);   multiplier m734(A[address][30],B[30][22],mul734);   multiplier m735(A[address][31],B[31][22],mul735);   
	multiplier m736(A[address][0],B[0][23],mul736);   multiplier m737(A[address][1],B[1][23],mul737);   multiplier m738(A[address][2],B[2][23],mul738);   multiplier m739(A[address][3],B[3][23],mul739);   multiplier m740(A[address][4],B[4][23],mul740);   multiplier m741(A[address][5],B[5][23],mul741);   multiplier m742(A[address][6],B[6][23],mul742);   multiplier m743(A[address][7],B[7][23],mul743);   multiplier m744(A[address][8],B[8][23],mul744);   multiplier m745(A[address][9],B[9][23],mul745);   multiplier m746(A[address][10],B[10][23],mul746);   multiplier m747(A[address][11],B[11][23],mul747);   multiplier m748(A[address][12],B[12][23],mul748);   multiplier m749(A[address][13],B[13][23],mul749);   multiplier m750(A[address][14],B[14][23],mul750);   multiplier m751(A[address][15],B[15][23],mul751);   multiplier m752(A[address][16],B[16][23],mul752);   multiplier m753(A[address][17],B[17][23],mul753);   multiplier m754(A[address][18],B[18][23],mul754);   multiplier m755(A[address][19],B[19][23],mul755);   multiplier m756(A[address][20],B[20][23],mul756);   multiplier m757(A[address][21],B[21][23],mul757);   multiplier m758(A[address][22],B[22][23],mul758);   multiplier m759(A[address][23],B[23][23],mul759);   multiplier m760(A[address][24],B[24][23],mul760);   multiplier m761(A[address][25],B[25][23],mul761);   multiplier m762(A[address][26],B[26][23],mul762);   multiplier m763(A[address][27],B[27][23],mul763);   multiplier m764(A[address][28],B[28][23],mul764);   multiplier m765(A[address][29],B[29][23],mul765);   multiplier m766(A[address][30],B[30][23],mul766);   multiplier m767(A[address][31],B[31][23],mul767);   
	multiplier m768(A[address][0],B[0][24],mul768);   multiplier m769(A[address][1],B[1][24],mul769);   multiplier m770(A[address][2],B[2][24],mul770);   multiplier m771(A[address][3],B[3][24],mul771);   multiplier m772(A[address][4],B[4][24],mul772);   multiplier m773(A[address][5],B[5][24],mul773);   multiplier m774(A[address][6],B[6][24],mul774);   multiplier m775(A[address][7],B[7][24],mul775);   multiplier m776(A[address][8],B[8][24],mul776);   multiplier m777(A[address][9],B[9][24],mul777);   multiplier m778(A[address][10],B[10][24],mul778);   multiplier m779(A[address][11],B[11][24],mul779);   multiplier m780(A[address][12],B[12][24],mul780);   multiplier m781(A[address][13],B[13][24],mul781);   multiplier m782(A[address][14],B[14][24],mul782);   multiplier m783(A[address][15],B[15][24],mul783);   multiplier m784(A[address][16],B[16][24],mul784);   multiplier m785(A[address][17],B[17][24],mul785);   multiplier m786(A[address][18],B[18][24],mul786);   multiplier m787(A[address][19],B[19][24],mul787);   multiplier m788(A[address][20],B[20][24],mul788);   multiplier m789(A[address][21],B[21][24],mul789);   multiplier m790(A[address][22],B[22][24],mul790);   multiplier m791(A[address][23],B[23][24],mul791);   multiplier m792(A[address][24],B[24][24],mul792);   multiplier m793(A[address][25],B[25][24],mul793);   multiplier m794(A[address][26],B[26][24],mul794);   multiplier m795(A[address][27],B[27][24],mul795);   multiplier m796(A[address][28],B[28][24],mul796);   multiplier m797(A[address][29],B[29][24],mul797);   multiplier m798(A[address][30],B[30][24],mul798);   multiplier m799(A[address][31],B[31][24],mul799);   
	multiplier m800(A[address][0],B[0][25],mul800);   multiplier m801(A[address][1],B[1][25],mul801);   multiplier m802(A[address][2],B[2][25],mul802);   multiplier m803(A[address][3],B[3][25],mul803);   multiplier m804(A[address][4],B[4][25],mul804);   multiplier m805(A[address][5],B[5][25],mul805);   multiplier m806(A[address][6],B[6][25],mul806);   multiplier m807(A[address][7],B[7][25],mul807);   multiplier m808(A[address][8],B[8][25],mul808);   multiplier m809(A[address][9],B[9][25],mul809);   multiplier m810(A[address][10],B[10][25],mul810);   multiplier m811(A[address][11],B[11][25],mul811);   multiplier m812(A[address][12],B[12][25],mul812);   multiplier m813(A[address][13],B[13][25],mul813);   multiplier m814(A[address][14],B[14][25],mul814);   multiplier m815(A[address][15],B[15][25],mul815);   multiplier m816(A[address][16],B[16][25],mul816);   multiplier m817(A[address][17],B[17][25],mul817);   multiplier m818(A[address][18],B[18][25],mul818);   multiplier m819(A[address][19],B[19][25],mul819);   multiplier m820(A[address][20],B[20][25],mul820);   multiplier m821(A[address][21],B[21][25],mul821);   multiplier m822(A[address][22],B[22][25],mul822);   multiplier m823(A[address][23],B[23][25],mul823);   multiplier m824(A[address][24],B[24][25],mul824);   multiplier m825(A[address][25],B[25][25],mul825);   multiplier m826(A[address][26],B[26][25],mul826);   multiplier m827(A[address][27],B[27][25],mul827);   multiplier m828(A[address][28],B[28][25],mul828);   multiplier m829(A[address][29],B[29][25],mul829);   multiplier m830(A[address][30],B[30][25],mul830);   multiplier m831(A[address][31],B[31][25],mul831);   
	multiplier m832(A[address][0],B[0][26],mul832);   multiplier m833(A[address][1],B[1][26],mul833);   multiplier m834(A[address][2],B[2][26],mul834);   multiplier m835(A[address][3],B[3][26],mul835);   multiplier m836(A[address][4],B[4][26],mul836);   multiplier m837(A[address][5],B[5][26],mul837);   multiplier m838(A[address][6],B[6][26],mul838);   multiplier m839(A[address][7],B[7][26],mul839);   multiplier m840(A[address][8],B[8][26],mul840);   multiplier m841(A[address][9],B[9][26],mul841);   multiplier m842(A[address][10],B[10][26],mul842);   multiplier m843(A[address][11],B[11][26],mul843);   multiplier m844(A[address][12],B[12][26],mul844);   multiplier m845(A[address][13],B[13][26],mul845);   multiplier m846(A[address][14],B[14][26],mul846);   multiplier m847(A[address][15],B[15][26],mul847);   multiplier m848(A[address][16],B[16][26],mul848);   multiplier m849(A[address][17],B[17][26],mul849);   multiplier m850(A[address][18],B[18][26],mul850);   multiplier m851(A[address][19],B[19][26],mul851);   multiplier m852(A[address][20],B[20][26],mul852);   multiplier m853(A[address][21],B[21][26],mul853);   multiplier m854(A[address][22],B[22][26],mul854);   multiplier m855(A[address][23],B[23][26],mul855);   multiplier m856(A[address][24],B[24][26],mul856);   multiplier m857(A[address][25],B[25][26],mul857);   multiplier m858(A[address][26],B[26][26],mul858);   multiplier m859(A[address][27],B[27][26],mul859);   multiplier m860(A[address][28],B[28][26],mul860);   multiplier m861(A[address][29],B[29][26],mul861);   multiplier m862(A[address][30],B[30][26],mul862);   multiplier m863(A[address][31],B[31][26],mul863);   
	multiplier m864(A[address][0],B[0][27],mul864);   multiplier m865(A[address][1],B[1][27],mul865);   multiplier m866(A[address][2],B[2][27],mul866);   multiplier m867(A[address][3],B[3][27],mul867);   multiplier m868(A[address][4],B[4][27],mul868);   multiplier m869(A[address][5],B[5][27],mul869);   multiplier m870(A[address][6],B[6][27],mul870);   multiplier m871(A[address][7],B[7][27],mul871);   multiplier m872(A[address][8],B[8][27],mul872);   multiplier m873(A[address][9],B[9][27],mul873);   multiplier m874(A[address][10],B[10][27],mul874);   multiplier m875(A[address][11],B[11][27],mul875);   multiplier m876(A[address][12],B[12][27],mul876);   multiplier m877(A[address][13],B[13][27],mul877);   multiplier m878(A[address][14],B[14][27],mul878);   multiplier m879(A[address][15],B[15][27],mul879);   multiplier m880(A[address][16],B[16][27],mul880);   multiplier m881(A[address][17],B[17][27],mul881);   multiplier m882(A[address][18],B[18][27],mul882);   multiplier m883(A[address][19],B[19][27],mul883);   multiplier m884(A[address][20],B[20][27],mul884);   multiplier m885(A[address][21],B[21][27],mul885);   multiplier m886(A[address][22],B[22][27],mul886);   multiplier m887(A[address][23],B[23][27],mul887);   multiplier m888(A[address][24],B[24][27],mul888);   multiplier m889(A[address][25],B[25][27],mul889);   multiplier m890(A[address][26],B[26][27],mul890);   multiplier m891(A[address][27],B[27][27],mul891);   multiplier m892(A[address][28],B[28][27],mul892);   multiplier m893(A[address][29],B[29][27],mul893);   multiplier m894(A[address][30],B[30][27],mul894);   multiplier m895(A[address][31],B[31][27],mul895);   
	multiplier m896(A[address][0],B[0][28],mul896);   multiplier m897(A[address][1],B[1][28],mul897);   multiplier m898(A[address][2],B[2][28],mul898);   multiplier m899(A[address][3],B[3][28],mul899);   multiplier m900(A[address][4],B[4][28],mul900);   multiplier m901(A[address][5],B[5][28],mul901);   multiplier m902(A[address][6],B[6][28],mul902);   multiplier m903(A[address][7],B[7][28],mul903);   multiplier m904(A[address][8],B[8][28],mul904);   multiplier m905(A[address][9],B[9][28],mul905);   multiplier m906(A[address][10],B[10][28],mul906);   multiplier m907(A[address][11],B[11][28],mul907);   multiplier m908(A[address][12],B[12][28],mul908);   multiplier m909(A[address][13],B[13][28],mul909);   multiplier m910(A[address][14],B[14][28],mul910);   multiplier m911(A[address][15],B[15][28],mul911);   multiplier m912(A[address][16],B[16][28],mul912);   multiplier m913(A[address][17],B[17][28],mul913);   multiplier m914(A[address][18],B[18][28],mul914);   multiplier m915(A[address][19],B[19][28],mul915);   multiplier m916(A[address][20],B[20][28],mul916);   multiplier m917(A[address][21],B[21][28],mul917);   multiplier m918(A[address][22],B[22][28],mul918);   multiplier m919(A[address][23],B[23][28],mul919);   multiplier m920(A[address][24],B[24][28],mul920);   multiplier m921(A[address][25],B[25][28],mul921);   multiplier m922(A[address][26],B[26][28],mul922);   multiplier m923(A[address][27],B[27][28],mul923);   multiplier m924(A[address][28],B[28][28],mul924);   multiplier m925(A[address][29],B[29][28],mul925);   multiplier m926(A[address][30],B[30][28],mul926);   multiplier m927(A[address][31],B[31][28],mul927);   
	multiplier m928(A[address][0],B[0][29],mul928);   multiplier m929(A[address][1],B[1][29],mul929);   multiplier m930(A[address][2],B[2][29],mul930);   multiplier m931(A[address][3],B[3][29],mul931);   multiplier m932(A[address][4],B[4][29],mul932);   multiplier m933(A[address][5],B[5][29],mul933);   multiplier m934(A[address][6],B[6][29],mul934);   multiplier m935(A[address][7],B[7][29],mul935);   multiplier m936(A[address][8],B[8][29],mul936);   multiplier m937(A[address][9],B[9][29],mul937);   multiplier m938(A[address][10],B[10][29],mul938);   multiplier m939(A[address][11],B[11][29],mul939);   multiplier m940(A[address][12],B[12][29],mul940);   multiplier m941(A[address][13],B[13][29],mul941);   multiplier m942(A[address][14],B[14][29],mul942);   multiplier m943(A[address][15],B[15][29],mul943);   multiplier m944(A[address][16],B[16][29],mul944);   multiplier m945(A[address][17],B[17][29],mul945);   multiplier m946(A[address][18],B[18][29],mul946);   multiplier m947(A[address][19],B[19][29],mul947);   multiplier m948(A[address][20],B[20][29],mul948);   multiplier m949(A[address][21],B[21][29],mul949);   multiplier m950(A[address][22],B[22][29],mul950);   multiplier m951(A[address][23],B[23][29],mul951);   multiplier m952(A[address][24],B[24][29],mul952);   multiplier m953(A[address][25],B[25][29],mul953);   multiplier m954(A[address][26],B[26][29],mul954);   multiplier m955(A[address][27],B[27][29],mul955);   multiplier m956(A[address][28],B[28][29],mul956);   multiplier m957(A[address][29],B[29][29],mul957);   multiplier m958(A[address][30],B[30][29],mul958);   multiplier m959(A[address][31],B[31][29],mul959);   
	multiplier m960(A[address][0],B[0][30],mul960);   multiplier m961(A[address][1],B[1][30],mul961);   multiplier m962(A[address][2],B[2][30],mul962);   multiplier m963(A[address][3],B[3][30],mul963);   multiplier m964(A[address][4],B[4][30],mul964);   multiplier m965(A[address][5],B[5][30],mul965);   multiplier m966(A[address][6],B[6][30],mul966);   multiplier m967(A[address][7],B[7][30],mul967);   multiplier m968(A[address][8],B[8][30],mul968);   multiplier m969(A[address][9],B[9][30],mul969);   multiplier m970(A[address][10],B[10][30],mul970);   multiplier m971(A[address][11],B[11][30],mul971);   multiplier m972(A[address][12],B[12][30],mul972);   multiplier m973(A[address][13],B[13][30],mul973);   multiplier m974(A[address][14],B[14][30],mul974);   multiplier m975(A[address][15],B[15][30],mul975);   multiplier m976(A[address][16],B[16][30],mul976);   multiplier m977(A[address][17],B[17][30],mul977);   multiplier m978(A[address][18],B[18][30],mul978);   multiplier m979(A[address][19],B[19][30],mul979);   multiplier m980(A[address][20],B[20][30],mul980);   multiplier m981(A[address][21],B[21][30],mul981);   multiplier m982(A[address][22],B[22][30],mul982);   multiplier m983(A[address][23],B[23][30],mul983);   multiplier m984(A[address][24],B[24][30],mul984);   multiplier m985(A[address][25],B[25][30],mul985);   multiplier m986(A[address][26],B[26][30],mul986);   multiplier m987(A[address][27],B[27][30],mul987);   multiplier m988(A[address][28],B[28][30],mul988);   multiplier m989(A[address][29],B[29][30],mul989);   multiplier m990(A[address][30],B[30][30],mul990);   multiplier m991(A[address][31],B[31][30],mul991);   
	multiplier m992(A[address][0],B[0][31],mul992);   multiplier m993(A[address][1],B[1][31],mul993);   multiplier m994(A[address][2],B[2][31],mul994);   multiplier m995(A[address][3],B[3][31],mul995);   multiplier m996(A[address][4],B[4][31],mul996);   multiplier m997(A[address][5],B[5][31],mul997);   multiplier m998(A[address][6],B[6][31],mul998);   multiplier m999(A[address][7],B[7][31],mul999);   multiplier m1000(A[address][8],B[8][31],mul1000);   multiplier m1001(A[address][9],B[9][31],mul1001);   multiplier m1002(A[address][10],B[10][31],mul1002);   multiplier m1003(A[address][11],B[11][31],mul1003);   multiplier m1004(A[address][12],B[12][31],mul1004);   multiplier m1005(A[address][13],B[13][31],mul1005);   multiplier m1006(A[address][14],B[14][31],mul1006);   multiplier m1007(A[address][15],B[15][31],mul1007);   multiplier m1008(A[address][16],B[16][31],mul1008);   multiplier m1009(A[address][17],B[17][31],mul1009);   multiplier m1010(A[address][18],B[18][31],mul1010);   multiplier m1011(A[address][19],B[19][31],mul1011);   multiplier m1012(A[address][20],B[20][31],mul1012);   multiplier m1013(A[address][21],B[21][31],mul1013);   multiplier m1014(A[address][22],B[22][31],mul1014);   multiplier m1015(A[address][23],B[23][31],mul1015);   multiplier m1016(A[address][24],B[24][31],mul1016);   multiplier m1017(A[address][25],B[25][31],mul1017);   multiplier m1018(A[address][26],B[26][31],mul1018);   multiplier m1019(A[address][27],B[27][31],mul1019);   multiplier m1020(A[address][28],B[28][31],mul1020);   multiplier m1021(A[address][29],B[29][31],mul1021);   multiplier m1022(A[address][30],B[30][31],mul1022);   multiplier m1023(A[address][31],B[31][31],mul1023);   

	
	adder a0(mul0,mul1,s0);   adder a1(s0,mul2,s1);   adder a2(s1,mul3,s2);   adder a3(s2,mul4,s3);   adder a4(s3,mul5,s4);   adder a5(s4,mul6,s5);   adder a6(s5,mul7,s6);   adder a7(s6,mul8,s7);   adder a8(s7,mul9,s8);   adder a9(s8,mul10,s9);   adder a10(s9,mul11,s10);   adder a11(s10,mul12,s11);   adder a12(s11,mul13,s12);   adder a13(s12,mul14,s13);   adder a14(s13,mul15,s14);   adder a15(s14,mul16,s15);   adder a16(s15,mul17,s16);   adder a17(s16,mul18,s17);   adder a18(s17,mul19,s18);   adder a19(s18,mul20,s19);   adder a20(s19,mul21,s20);   adder a21(s20,mul22,s21);   adder a22(s21,mul23,s22);   adder a23(s22,mul24,s23);   adder a24(s23,mul25,s24);   adder a25(s24,mul26,s25);   adder a26(s25,mul27,s26);   adder a27(s26,mul28,s27);   adder a28(s27,mul29,s28);   adder a29(s28,mul30,s29);   adder a30(s29,mul31,s30);   
	adder a32(mul32,mul33,s31);   adder a33(s31,mul34,s32);   adder a34(s32,mul35,s33);   adder a35(s33,mul36,s34);   adder a36(s34,mul37,s35);   adder a37(s35,mul38,s36);   adder a38(s36,mul39,s37);   adder a39(s37,mul40,s38);   adder a40(s38,mul41,s39);   adder a41(s39,mul42,s40);   adder a42(s40,mul43,s41);   adder a43(s41,mul44,s42);   adder a44(s42,mul45,s43);   adder a45(s43,mul46,s44);   adder a46(s44,mul47,s45);   adder a47(s45,mul48,s46);   adder a48(s46,mul49,s47);   adder a49(s47,mul50,s48);   adder a50(s48,mul51,s49);   adder a51(s49,mul52,s50);   adder a52(s50,mul53,s51);   adder a53(s51,mul54,s52);   adder a54(s52,mul55,s53);   adder a55(s53,mul56,s54);   adder a56(s54,mul57,s55);   adder a57(s55,mul58,s56);   adder a58(s56,mul59,s57);   adder a59(s57,mul60,s58);   adder a60(s58,mul61,s59);   adder a61(s59,mul62,s60);   adder a62(s60,mul63,s61);
   adder a64(mul64,mul65,s62);   adder a65(s62,mul66,s63);   adder a66(s63,mul67,s64);   adder a67(s64,mul68,s65);   adder a68(s65,mul69,s66);   adder a69(s66,mul70,s67);   adder a70(s67,mul71,s68);   adder a71(s68,mul72,s69);   adder a72(s69,mul73,s70);   adder a73(s70,mul74,s71);   adder a74(s71,mul75,s72);   adder a75(s72,mul76,s73);   adder a76(s73,mul77,s74);   adder a77(s74,mul78,s75);   adder a78(s75,mul79,s76);   adder a79(s76,mul80,s77);   adder a80(s77,mul81,s78);   adder a81(s78,mul82,s79);   adder a82(s79,mul83,s80);   adder a83(s80,mul84,s81);   adder a84(s81,mul85,s82);   adder a85(s82,mul86,s83);   adder a86(s83,mul87,s84);   adder a87(s84,mul88,s85);   adder a88(s85,mul89,s86);   adder a89(s86,mul90,s87);   adder a90(s87,mul91,s88);   adder a91(s88,mul92,s89);   adder a92(s89,mul93,s90);   adder a93(s90,mul94,s91);   adder a94(s91,mul95,s92);   
	adder a96(mul96,mul97,s93);   adder a97(s93,mul98,s94);   adder a98(s94,mul99,s95);   adder a99(s95,mul100,s96);   adder a100(s96,mul101,s97);   adder a101(s97,mul102,s98);   adder a102(s98,mul103,s99);   adder a103(s99,mul104,s100);   adder a104(s100,mul105,s101);   adder a105(s101,mul106,s102);   adder a106(s102,mul107,s103);   adder a107(s103,mul108,s104);   adder a108(s104,mul109,s105);   adder a109(s105,mul110,s106);   adder a110(s106,mul111,s107);   adder a111(s107,mul112,s108);   adder a112(s108,mul113,s109);   adder a113(s109,mul114,s110);   adder a114(s110,mul115,s111);   adder a115(s111,mul116,s112);   adder a116(s112,mul117,s113);   adder a117(s113,mul118,s114);   adder a118(s114,mul119,s115);   adder a119(s115,mul120,s116);   adder a120(s116,mul121,s117);   adder a121(s117,mul122,s118);   adder a122(s118,mul123,s119);   adder a123(s119,mul124,s120);   adder a124(s120,mul125,s121);   adder a125(s121,mul126,s122);   adder a126(s122,mul127,s123);   
	adder a128(mul128,mul129,s124);   adder a129(s124,mul130,s125);   adder a130(s125,mul131,s126);   adder a131(s126,mul132,s127);   adder a132(s127,mul133,s128);   adder a133(s128,mul134,s129);   adder a134(s129,mul135,s130);   adder a135(s130,mul136,s131);   adder a136(s131,mul137,s132);   adder a137(s132,mul138,s133);   adder a138(s133,mul139,s134);   adder a139(s134,mul140,s135);   adder a140(s135,mul141,s136);   adder a141(s136,mul142,s137);   adder a142(s137,mul143,s138);   adder a143(s138,mul144,s139);   adder a144(s139,mul145,s140);   adder a145(s140,mul146,s141);   adder a146(s141,mul147,s142);   adder a147(s142,mul148,s143);   adder a148(s143,mul149,s144);   adder a149(s144,mul150,s145);   adder a150(s145,mul151,s146);   adder a151(s146,mul152,s147);   adder a152(s147,mul153,s148);   adder a153(s148,mul154,s149);   adder a154(s149,mul155,s150);   adder a155(s150,mul156,s151);   adder a156(s151,mul157,s152);   adder a157(s152,mul158,s153);   adder a158(s153,mul159,s154);   
	adder a160(mul160,mul161,s155);   adder a161(s155,mul162,s156);   adder a162(s156,mul163,s157);   adder a163(s157,mul164,s158);   adder a164(s158,mul165,s159);   adder a165(s159,mul166,s160);   adder a166(s160,mul167,s161);   adder a167(s161,mul168,s162);   adder a168(s162,mul169,s163);   adder a169(s163,mul170,s164);   adder a170(s164,mul171,s165);   adder a171(s165,mul172,s166);   adder a172(s166,mul173,s167);   adder a173(s167,mul174,s168);   adder a174(s168,mul175,s169);   adder a175(s169,mul176,s170);   adder a176(s170,mul177,s171);   adder a177(s171,mul178,s172);   adder a178(s172,mul179,s173);   adder a179(s173,mul180,s174);   adder a180(s174,mul181,s175);   adder a181(s175,mul182,s176);   adder a182(s176,mul183,s177);   adder a183(s177,mul184,s178);   adder a184(s178,mul185,s179);   adder a185(s179,mul186,s180);   adder a186(s180,mul187,s181);   adder a187(s181,mul188,s182);   adder a188(s182,mul189,s183);   adder a189(s183,mul190,s184);   adder a190(s184,mul191,s185);   
	adder a192(mul192,mul193,s186);   adder a193(s186,mul194,s187);   adder a194(s187,mul195,s188);   adder a195(s188,mul196,s189);   adder a196(s189,mul197,s190);   adder a197(s190,mul198,s191);   adder a198(s191,mul199,s192);   adder a199(s192,mul200,s193);   adder a200(s193,mul201,s194);   adder a201(s194,mul202,s195);   adder a202(s195,mul203,s196);   adder a203(s196,mul204,s197);   adder a204(s197,mul205,s198);   adder a205(s198,mul206,s199);   adder a206(s199,mul207,s200);   adder a207(s200,mul208,s201);   adder a208(s201,mul209,s202);   adder a209(s202,mul210,s203);   adder a210(s203,mul211,s204);   adder a211(s204,mul212,s205);   adder a212(s205,mul213,s206);   adder a213(s206,mul214,s207);   adder a214(s207,mul215,s208);   adder a215(s208,mul216,s209);   adder a216(s209,mul217,s210);   adder a217(s210,mul218,s211);   adder a218(s211,mul219,s212);   adder a219(s212,mul220,s213);   adder a220(s213,mul221,s214);   adder a221(s214,mul222,s215);   adder a222(s215,mul223,s216);   
	adder a224(mul224,mul225,s217);   adder a225(s217,mul226,s218);   adder a226(s218,mul227,s219);   adder a227(s219,mul228,s220);   adder a228(s220,mul229,s221);   adder a229(s221,mul230,s222);   adder a230(s222,mul231,s223);   adder a231(s223,mul232,s224);   adder a232(s224,mul233,s225);   adder a233(s225,mul234,s226);   adder a234(s226,mul235,s227);   adder a235(s227,mul236,s228);   adder a236(s228,mul237,s229);   adder a237(s229,mul238,s230);   adder a238(s230,mul239,s231);   adder a239(s231,mul240,s232);   adder a240(s232,mul241,s233);   adder a241(s233,mul242,s234);   adder a242(s234,mul243,s235);   adder a243(s235,mul244,s236);   adder a244(s236,mul245,s237);   adder a245(s237,mul246,s238);   adder a246(s238,mul247,s239);   adder a247(s239,mul248,s240);   adder a248(s240,mul249,s241);   adder a249(s241,mul250,s242);   adder a250(s242,mul251,s243);   adder a251(s243,mul252,s244);   adder a252(s244,mul253,s245);   adder a253(s245,mul254,s246);   adder a254(s246,mul255,s247);   
	adder a256(mul256,mul257,s248);   adder a257(s248,mul258,s249);   adder a258(s249,mul259,s250);   adder a259(s250,mul260,s251);   adder a260(s251,mul261,s252);   adder a261(s252,mul262,s253);   adder a262(s253,mul263,s254);   adder a263(s254,mul264,s255);   adder a264(s255,mul265,s256);   adder a265(s256,mul266,s257);   adder a266(s257,mul267,s258);   adder a267(s258,mul268,s259);   adder a268(s259,mul269,s260);   adder a269(s260,mul270,s261);   adder a270(s261,mul271,s262);   adder a271(s262,mul272,s263);   adder a272(s263,mul273,s264);   adder a273(s264,mul274,s265);   adder a274(s265,mul275,s266);   adder a275(s266,mul276,s267);   adder a276(s267,mul277,s268);   adder a277(s268,mul278,s269);   adder a278(s269,mul279,s270);   adder a279(s270,mul280,s271);   adder a280(s271,mul281,s272);   adder a281(s272,mul282,s273);   adder a282(s273,mul283,s274);   adder a283(s274,mul284,s275);   adder a284(s275,mul285,s276);   adder a285(s276,mul286,s277);   adder a286(s277,mul287,s278);   
	adder a288(mul288,mul289,s279);   adder a289(s279,mul290,s280);   adder a290(s280,mul291,s281);   adder a291(s281,mul292,s282);   adder a292(s282,mul293,s283);   adder a293(s283,mul294,s284);   adder a294(s284,mul295,s285);   adder a295(s285,mul296,s286);   adder a296(s286,mul297,s287);   adder a297(s287,mul298,s288);   adder a298(s288,mul299,s289);   adder a299(s289,mul300,s290);   adder a300(s290,mul301,s291);   adder a301(s291,mul302,s292);   adder a302(s292,mul303,s293);   adder a303(s293,mul304,s294);   adder a304(s294,mul305,s295);   adder a305(s295,mul306,s296);   adder a306(s296,mul307,s297);   adder a307(s297,mul308,s298);   adder a308(s298,mul309,s299);   adder a309(s299,mul310,s300);   adder a310(s300,mul311,s301);   adder a311(s301,mul312,s302);   adder a312(s302,mul313,s303);   adder a313(s303,mul314,s304);   adder a314(s304,mul315,s305);   adder a315(s305,mul316,s306);   adder a316(s306,mul317,s307);   adder a317(s307,mul318,s308);   adder a318(s308,mul319,s309);   
	adder a320(mul320,mul321,s310);   adder a321(s310,mul322,s311);   adder a322(s311,mul323,s312);   adder a323(s312,mul324,s313);   adder a324(s313,mul325,s314);   adder a325(s314,mul326,s315);   adder a326(s315,mul327,s316);   adder a327(s316,mul328,s317);   adder a328(s317,mul329,s318);   adder a329(s318,mul330,s319);   adder a330(s319,mul331,s320);   adder a331(s320,mul332,s321);   adder a332(s321,mul333,s322);   adder a333(s322,mul334,s323);   adder a334(s323,mul335,s324);   adder a335(s324,mul336,s325);   adder a336(s325,mul337,s326);   adder a337(s326,mul338,s327);   adder a338(s327,mul339,s328);   adder a339(s328,mul340,s329);   adder a340(s329,mul341,s330);   adder a341(s330,mul342,s331);   adder a342(s331,mul343,s332);   adder a343(s332,mul344,s333);   adder a344(s333,mul345,s334);   adder a345(s334,mul346,s335);   adder a346(s335,mul347,s336);   adder a347(s336,mul348,s337);   adder a348(s337,mul349,s338);   adder a349(s338,mul350,s339);   adder a350(s339,mul351,s340);   
	adder a352(mul352,mul353,s341);   adder a353(s341,mul354,s342);   adder a354(s342,mul355,s343);   adder a355(s343,mul356,s344);   adder a356(s344,mul357,s345);   adder a357(s345,mul358,s346);   adder a358(s346,mul359,s347);   adder a359(s347,mul360,s348);   adder a360(s348,mul361,s349);   adder a361(s349,mul362,s350);   adder a362(s350,mul363,s351);   adder a363(s351,mul364,s352);   adder a364(s352,mul365,s353);   adder a365(s353,mul366,s354);   adder a366(s354,mul367,s355);   adder a367(s355,mul368,s356);   adder a368(s356,mul369,s357);   adder a369(s357,mul370,s358);   adder a370(s358,mul371,s359);   adder a371(s359,mul372,s360);   adder a372(s360,mul373,s361);   adder a373(s361,mul374,s362);   adder a374(s362,mul375,s363);   adder a375(s363,mul376,s364);   adder a376(s364,mul377,s365);   adder a377(s365,mul378,s366);   adder a378(s366,mul379,s367);   adder a379(s367,mul380,s368);   adder a380(s368,mul381,s369);   adder a381(s369,mul382,s370);   adder a382(s370,mul383,s371);   
	adder a384(mul384,mul385,s372);   adder a385(s372,mul386,s373);   adder a386(s373,mul387,s374);   adder a387(s374,mul388,s375);   adder a388(s375,mul389,s376);   adder a389(s376,mul390,s377);   adder a390(s377,mul391,s378);   adder a391(s378,mul392,s379);   adder a392(s379,mul393,s380);   adder a393(s380,mul394,s381);   adder a394(s381,mul395,s382);   adder a395(s382,mul396,s383);   adder a396(s383,mul397,s384);   adder a397(s384,mul398,s385);   adder a398(s385,mul399,s386);   adder a399(s386,mul400,s387);   adder a400(s387,mul401,s388);   adder a401(s388,mul402,s389);   adder a402(s389,mul403,s390);   adder a403(s390,mul404,s391);   adder a404(s391,mul405,s392);   adder a405(s392,mul406,s393);   adder a406(s393,mul407,s394);   adder a407(s394,mul408,s395);   adder a408(s395,mul409,s396);   adder a409(s396,mul410,s397);   adder a410(s397,mul411,s398);   adder a411(s398,mul412,s399);   adder a412(s399,mul413,s400);   adder a413(s400,mul414,s401);   adder a414(s401,mul415,s402);   
	adder a416(mul416,mul417,s403);   adder a417(s403,mul418,s404);   adder a418(s404,mul419,s405);   adder a419(s405,mul420,s406);   adder a420(s406,mul421,s407);   adder a421(s407,mul422,s408);   adder a422(s408,mul423,s409);   adder a423(s409,mul424,s410);   adder a424(s410,mul425,s411);   adder a425(s411,mul426,s412);   adder a426(s412,mul427,s413);   adder a427(s413,mul428,s414);   adder a428(s414,mul429,s415);   adder a429(s415,mul430,s416);   adder a430(s416,mul431,s417);   adder a431(s417,mul432,s418);   adder a432(s418,mul433,s419);   adder a433(s419,mul434,s420);   adder a434(s420,mul435,s421);   adder a435(s421,mul436,s422);   adder a436(s422,mul437,s423);   adder a437(s423,mul438,s424);   adder a438(s424,mul439,s425);   adder a439(s425,mul440,s426);   adder a440(s426,mul441,s427);   adder a441(s427,mul442,s428);   adder a442(s428,mul443,s429);   adder a443(s429,mul444,s430);   adder a444(s430,mul445,s431);   adder a445(s431,mul446,s432);   adder a446(s432,mul447,s433);   
	adder a448(mul448,mul449,s434);   adder a449(s434,mul450,s435);   adder a450(s435,mul451,s436);   adder a451(s436,mul452,s437);   adder a452(s437,mul453,s438);   adder a453(s438,mul454,s439);   adder a454(s439,mul455,s440);   adder a455(s440,mul456,s441);   adder a456(s441,mul457,s442);   adder a457(s442,mul458,s443);   adder a458(s443,mul459,s444);   adder a459(s444,mul460,s445);   adder a460(s445,mul461,s446);   adder a461(s446,mul462,s447);   adder a462(s447,mul463,s448);   adder a463(s448,mul464,s449);   adder a464(s449,mul465,s450);   adder a465(s450,mul466,s451);   adder a466(s451,mul467,s452);   adder a467(s452,mul468,s453);   adder a468(s453,mul469,s454);   adder a469(s454,mul470,s455);   adder a470(s455,mul471,s456);   adder a471(s456,mul472,s457);   adder a472(s457,mul473,s458);   adder a473(s458,mul474,s459);   adder a474(s459,mul475,s460);   adder a475(s460,mul476,s461);   adder a476(s461,mul477,s462);   adder a477(s462,mul478,s463);   adder a478(s463,mul479,s464);   
	adder a480(mul480,mul481,s465);   adder a481(s465,mul482,s466);   adder a482(s466,mul483,s467);   adder a483(s467,mul484,s468);   adder a484(s468,mul485,s469);   adder a485(s469,mul486,s470);   adder a486(s470,mul487,s471);   adder a487(s471,mul488,s472);   adder a488(s472,mul489,s473);   adder a489(s473,mul490,s474);   adder a490(s474,mul491,s475);   adder a491(s475,mul492,s476);   adder a492(s476,mul493,s477);   adder a493(s477,mul494,s478);   adder a494(s478,mul495,s479);   adder a495(s479,mul496,s480);   adder a496(s480,mul497,s481);   adder a497(s481,mul498,s482);   adder a498(s482,mul499,s483);   adder a499(s483,mul500,s484);   adder a500(s484,mul501,s485);   adder a501(s485,mul502,s486);   adder a502(s486,mul503,s487);   adder a503(s487,mul504,s488);   adder a504(s488,mul505,s489);   adder a505(s489,mul506,s490);   adder a506(s490,mul507,s491);   adder a507(s491,mul508,s492);   adder a508(s492,mul509,s493);   adder a509(s493,mul510,s494);   adder a510(s494,mul511,s495);   
	adder a512(mul512,mul513,s496);   adder a513(s496,mul514,s497);   adder a514(s497,mul515,s498);   adder a515(s498,mul516,s499);   adder a516(s499,mul517,s500);   adder a517(s500,mul518,s501);   adder a518(s501,mul519,s502);   adder a519(s502,mul520,s503);   adder a520(s503,mul521,s504);   adder a521(s504,mul522,s505);   adder a522(s505,mul523,s506);   adder a523(s506,mul524,s507);   adder a524(s507,mul525,s508);   adder a525(s508,mul526,s509);   adder a526(s509,mul527,s510);   adder a527(s510,mul528,s511);   adder a528(s511,mul529,s512);   adder a529(s512,mul530,s513);   adder a530(s513,mul531,s514);   adder a531(s514,mul532,s515);   adder a532(s515,mul533,s516);   adder a533(s516,mul534,s517);   adder a534(s517,mul535,s518);   adder a535(s518,mul536,s519);   adder a536(s519,mul537,s520);   adder a537(s520,mul538,s521);   adder a538(s521,mul539,s522);   adder a539(s522,mul540,s523);   adder a540(s523,mul541,s524);   adder a541(s524,mul542,s525);   adder a542(s525,mul543,s526);   
	adder a544(mul544,mul545,s527);   adder a545(s527,mul546,s528);   adder a546(s528,mul547,s529);   adder a547(s529,mul548,s530);   adder a548(s530,mul549,s531);   adder a549(s531,mul550,s532);   adder a550(s532,mul551,s533);   adder a551(s533,mul552,s534);   adder a552(s534,mul553,s535);   adder a553(s535,mul554,s536);   adder a554(s536,mul555,s537);   adder a555(s537,mul556,s538);   adder a556(s538,mul557,s539);   adder a557(s539,mul558,s540);   adder a558(s540,mul559,s541);   adder a559(s541,mul560,s542);   adder a560(s542,mul561,s543);   adder a561(s543,mul562,s544);   adder a562(s544,mul563,s545);   adder a563(s545,mul564,s546);   adder a564(s546,mul565,s547);   adder a565(s547,mul566,s548);   adder a566(s548,mul567,s549);   adder a567(s549,mul568,s550);   adder a568(s550,mul569,s551);   adder a569(s551,mul570,s552);   adder a570(s552,mul571,s553);   adder a571(s553,mul572,s554);   adder a572(s554,mul573,s555);   adder a573(s555,mul574,s556);   adder a574(s556,mul575,s557);   
	adder a576(mul576,mul577,s558);   adder a577(s558,mul578,s559);   adder a578(s559,mul579,s560);   adder a579(s560,mul580,s561);   adder a580(s561,mul581,s562);   adder a581(s562,mul582,s563);   adder a582(s563,mul583,s564);   adder a583(s564,mul584,s565);   adder a584(s565,mul585,s566);   adder a585(s566,mul586,s567);   adder a586(s567,mul587,s568);   adder a587(s568,mul588,s569);   adder a588(s569,mul589,s570);   adder a589(s570,mul590,s571);   adder a590(s571,mul591,s572);   adder a591(s572,mul592,s573);   adder a592(s573,mul593,s574);   adder a593(s574,mul594,s575);   adder a594(s575,mul595,s576);   adder a595(s576,mul596,s577);   adder a596(s577,mul597,s578);   adder a597(s578,mul598,s579);   adder a598(s579,mul599,s580);   adder a599(s580,mul600,s581);   adder a600(s581,mul601,s582);   adder a601(s582,mul602,s583);   adder a602(s583,mul603,s584);   adder a603(s584,mul604,s585);   adder a604(s585,mul605,s586);   adder a605(s586,mul606,s587);   adder a606(s587,mul607,s588);   
	adder a608(mul608,mul609,s589);   adder a609(s589,mul610,s590);   adder a610(s590,mul611,s591);   adder a611(s591,mul612,s592);   adder a612(s592,mul613,s593);   adder a613(s593,mul614,s594);   adder a614(s594,mul615,s595);   adder a615(s595,mul616,s596);   adder a616(s596,mul617,s597);   adder a617(s597,mul618,s598);   adder a618(s598,mul619,s599);   adder a619(s599,mul620,s600);   adder a620(s600,mul621,s601);   adder a621(s601,mul622,s602);   adder a622(s602,mul623,s603);   adder a623(s603,mul624,s604);   adder a624(s604,mul625,s605);   adder a625(s605,mul626,s606);   adder a626(s606,mul627,s607);   adder a627(s607,mul628,s608);   adder a628(s608,mul629,s609);   adder a629(s609,mul630,s610);   adder a630(s610,mul631,s611);   adder a631(s611,mul632,s612);   adder a632(s612,mul633,s613);   adder a633(s613,mul634,s614);   adder a634(s614,mul635,s615);   adder a635(s615,mul636,s616);   adder a636(s616,mul637,s617);   adder a637(s617,mul638,s618);   adder a638(s618,mul639,s619);   
	adder a640(mul640,mul641,s620);   adder a641(s620,mul642,s621);   adder a642(s621,mul643,s622);   adder a643(s622,mul644,s623);   adder a644(s623,mul645,s624);   adder a645(s624,mul646,s625);   adder a646(s625,mul647,s626);   adder a647(s626,mul648,s627);   adder a648(s627,mul649,s628);   adder a649(s628,mul650,s629);   adder a650(s629,mul651,s630);   adder a651(s630,mul652,s631);   adder a652(s631,mul653,s632);   adder a653(s632,mul654,s633);   adder a654(s633,mul655,s634);   adder a655(s634,mul656,s635);   adder a656(s635,mul657,s636);   adder a657(s636,mul658,s637);   adder a658(s637,mul659,s638);   adder a659(s638,mul660,s639);   adder a660(s639,mul661,s640);   adder a661(s640,mul662,s641);   adder a662(s641,mul663,s642);   adder a663(s642,mul664,s643);   adder a664(s643,mul665,s644);   adder a665(s644,mul666,s645);   adder a666(s645,mul667,s646);   adder a667(s646,mul668,s647);   adder a668(s647,mul669,s648);   adder a669(s648,mul670,s649);   adder a670(s649,mul671,s650);   
	adder a672(mul672,mul673,s651);   adder a673(s651,mul674,s652);   adder a674(s652,mul675,s653);   adder a675(s653,mul676,s654);   adder a676(s654,mul677,s655);   adder a677(s655,mul678,s656);   adder a678(s656,mul679,s657);   adder a679(s657,mul680,s658);   adder a680(s658,mul681,s659);   adder a681(s659,mul682,s660);   adder a682(s660,mul683,s661);   adder a683(s661,mul684,s662);   adder a684(s662,mul685,s663);   adder a685(s663,mul686,s664);   adder a686(s664,mul687,s665);   adder a687(s665,mul688,s666);   adder a688(s666,mul689,s667);   adder a689(s667,mul690,s668);   adder a690(s668,mul691,s669);   adder a691(s669,mul692,s670);   adder a692(s670,mul693,s671);   adder a693(s671,mul694,s672);   adder a694(s672,mul695,s673);   adder a695(s673,mul696,s674);   adder a696(s674,mul697,s675);   adder a697(s675,mul698,s676);   adder a698(s676,mul699,s677);   adder a699(s677,mul700,s678);   adder a700(s678,mul701,s679);   adder a701(s679,mul702,s680);   adder a702(s680,mul703,s681);   
	adder a704(mul704,mul705,s682);   adder a705(s682,mul706,s683);   adder a706(s683,mul707,s684);   adder a707(s684,mul708,s685);   adder a708(s685,mul709,s686);   adder a709(s686,mul710,s687);   adder a710(s687,mul711,s688);   adder a711(s688,mul712,s689);   adder a712(s689,mul713,s690);   adder a713(s690,mul714,s691);   adder a714(s691,mul715,s692);   adder a715(s692,mul716,s693);   adder a716(s693,mul717,s694);   adder a717(s694,mul718,s695);   adder a718(s695,mul719,s696);   adder a719(s696,mul720,s697);   adder a720(s697,mul721,s698);   adder a721(s698,mul722,s699);   adder a722(s699,mul723,s700);   adder a723(s700,mul724,s701);   adder a724(s701,mul725,s702);   adder a725(s702,mul726,s703);   adder a726(s703,mul727,s704);   adder a727(s704,mul728,s705);   adder a728(s705,mul729,s706);   adder a729(s706,mul730,s707);   adder a730(s707,mul731,s708);   adder a731(s708,mul732,s709);   adder a732(s709,mul733,s710);   adder a733(s710,mul734,s711);   adder a734(s711,mul735,s712);   
	adder a736(mul736,mul737,s713);   adder a737(s713,mul738,s714);   adder a738(s714,mul739,s715);   adder a739(s715,mul740,s716);   adder a740(s716,mul741,s717);   adder a741(s717,mul742,s718);   adder a742(s718,mul743,s719);   adder a743(s719,mul744,s720);   adder a744(s720,mul745,s721);   adder a745(s721,mul746,s722);   adder a746(s722,mul747,s723);   adder a747(s723,mul748,s724);   adder a748(s724,mul749,s725);   adder a749(s725,mul750,s726);   adder a750(s726,mul751,s727);   adder a751(s727,mul752,s728);   adder a752(s728,mul753,s729);   adder a753(s729,mul754,s730);   adder a754(s730,mul755,s731);   adder a755(s731,mul756,s732);   adder a756(s732,mul757,s733);   adder a757(s733,mul758,s734);   adder a758(s734,mul759,s735);   adder a759(s735,mul760,s736);   adder a760(s736,mul761,s737);   adder a761(s737,mul762,s738);   adder a762(s738,mul763,s739);   adder a763(s739,mul764,s740);   adder a764(s740,mul765,s741);   adder a765(s741,mul766,s742);   adder a766(s742,mul767,s743);   
	adder a768(mul768,mul769,s744);   adder a769(s744,mul770,s745);   adder a770(s745,mul771,s746);   adder a771(s746,mul772,s747);   adder a772(s747,mul773,s748);   adder a773(s748,mul774,s749);   adder a774(s749,mul775,s750);   adder a775(s750,mul776,s751);   adder a776(s751,mul777,s752);   adder a777(s752,mul778,s753);   adder a778(s753,mul779,s754);   adder a779(s754,mul780,s755);   adder a780(s755,mul781,s756);   adder a781(s756,mul782,s757);   adder a782(s757,mul783,s758);   adder a783(s758,mul784,s759);   adder a784(s759,mul785,s760);   adder a785(s760,mul786,s761);   adder a786(s761,mul787,s762);   adder a787(s762,mul788,s763);   adder a788(s763,mul789,s764);   adder a789(s764,mul790,s765);   adder a790(s765,mul791,s766);   adder a791(s766,mul792,s767);   adder a792(s767,mul793,s768);   adder a793(s768,mul794,s769);   adder a794(s769,mul795,s770);   adder a795(s770,mul796,s771);   adder a796(s771,mul797,s772);   adder a797(s772,mul798,s773);   adder a798(s773,mul799,s774);   
	adder a800(mul800,mul801,s775);   adder a801(s775,mul802,s776);   adder a802(s776,mul803,s777);   adder a803(s777,mul804,s778);   adder a804(s778,mul805,s779);   adder a805(s779,mul806,s780);   adder a806(s780,mul807,s781);   adder a807(s781,mul808,s782);   adder a808(s782,mul809,s783);   adder a809(s783,mul810,s784);   adder a810(s784,mul811,s785);   adder a811(s785,mul812,s786);   adder a812(s786,mul813,s787);   adder a813(s787,mul814,s788);   adder a814(s788,mul815,s789);   adder a815(s789,mul816,s790);   adder a816(s790,mul817,s791);   adder a817(s791,mul818,s792);   adder a818(s792,mul819,s793);   adder a819(s793,mul820,s794);   adder a820(s794,mul821,s795);   adder a821(s795,mul822,s796);   adder a822(s796,mul823,s797);   adder a823(s797,mul824,s798);   adder a824(s798,mul825,s799);   adder a825(s799,mul826,s800);   adder a826(s800,mul827,s801);   adder a827(s801,mul828,s802);   adder a828(s802,mul829,s803);   adder a829(s803,mul830,s804);   adder a830(s804,mul831,s805);   
	adder a832(mul832,mul833,s806);   adder a833(s806,mul834,s807);   adder a834(s807,mul835,s808);   adder a835(s808,mul836,s809);   adder a836(s809,mul837,s810);   adder a837(s810,mul838,s811);   adder a838(s811,mul839,s812);   adder a839(s812,mul840,s813);   adder a840(s813,mul841,s814);   adder a841(s814,mul842,s815);   adder a842(s815,mul843,s816);   adder a843(s816,mul844,s817);   adder a844(s817,mul845,s818);   adder a845(s818,mul846,s819);   adder a846(s819,mul847,s820);   adder a847(s820,mul848,s821);   adder a848(s821,mul849,s822);   adder a849(s822,mul850,s823);   adder a850(s823,mul851,s824);   adder a851(s824,mul852,s825);   adder a852(s825,mul853,s826);   adder a853(s826,mul854,s827);   adder a854(s827,mul855,s828);   adder a855(s828,mul856,s829);   adder a856(s829,mul857,s830);   adder a857(s830,mul858,s831);   adder a858(s831,mul859,s832);   adder a859(s832,mul860,s833);   adder a860(s833,mul861,s834);   adder a861(s834,mul862,s835);   adder a862(s835,mul863,s836);   
	adder a864(mul864,mul865,s837);   adder a865(s837,mul866,s838);   adder a866(s838,mul867,s839);   adder a867(s839,mul868,s840);   adder a868(s840,mul869,s841);   adder a869(s841,mul870,s842);   adder a870(s842,mul871,s843);   adder a871(s843,mul872,s844);   adder a872(s844,mul873,s845);   adder a873(s845,mul874,s846);   adder a874(s846,mul875,s847);   adder a875(s847,mul876,s848);   adder a876(s848,mul877,s849);   adder a877(s849,mul878,s850);   adder a878(s850,mul879,s851);   adder a879(s851,mul880,s852);   adder a880(s852,mul881,s853);   adder a881(s853,mul882,s854);   adder a882(s854,mul883,s855);   adder a883(s855,mul884,s856);   adder a884(s856,mul885,s857);   adder a885(s857,mul886,s858);   adder a886(s858,mul887,s859);   adder a887(s859,mul888,s860);   adder a888(s860,mul889,s861);   adder a889(s861,mul890,s862);   adder a890(s862,mul891,s863);   adder a891(s863,mul892,s864);   adder a892(s864,mul893,s865);   adder a893(s865,mul894,s866);   adder a894(s866,mul895,s867);   
	adder a896(mul896,mul897,s868);   adder a897(s868,mul898,s869);   adder a898(s869,mul899,s870);   adder a899(s870,mul900,s871);   adder a900(s871,mul901,s872);   adder a901(s872,mul902,s873);   adder a902(s873,mul903,s874);   adder a903(s874,mul904,s875);   adder a904(s875,mul905,s876);   adder a905(s876,mul906,s877);   adder a906(s877,mul907,s878);   adder a907(s878,mul908,s879);   adder a908(s879,mul909,s880);   adder a909(s880,mul910,s881);   adder a910(s881,mul911,s882);   adder a911(s882,mul912,s883);   adder a912(s883,mul913,s884);   adder a913(s884,mul914,s885);   adder a914(s885,mul915,s886);   adder a915(s886,mul916,s887);   adder a916(s887,mul917,s888);   adder a917(s888,mul918,s889);   adder a918(s889,mul919,s890);   adder a919(s890,mul920,s891);   adder a920(s891,mul921,s892);   adder a921(s892,mul922,s893);   adder a922(s893,mul923,s894);   adder a923(s894,mul924,s895);   adder a924(s895,mul925,s896);   adder a925(s896,mul926,s897);   adder a926(s897,mul927,s898);   
	adder a928(mul928,mul929,s899);   adder a929(s899,mul930,s900);   adder a930(s900,mul931,s901);   adder a931(s901,mul932,s902);   adder a932(s902,mul933,s903);   adder a933(s903,mul934,s904);   adder a934(s904,mul935,s905);   adder a935(s905,mul936,s906);   adder a936(s906,mul937,s907);   adder a937(s907,mul938,s908);   adder a938(s908,mul939,s909);   adder a939(s909,mul940,s910);   adder a940(s910,mul941,s911);   adder a941(s911,mul942,s912);   adder a942(s912,mul943,s913);   adder a943(s913,mul944,s914);   adder a944(s914,mul945,s915);   adder a945(s915,mul946,s916);   adder a946(s916,mul947,s917);   adder a947(s917,mul948,s918);   adder a948(s918,mul949,s919);   adder a949(s919,mul950,s920);   adder a950(s920,mul951,s921);   adder a951(s921,mul952,s922);   adder a952(s922,mul953,s923);   adder a953(s923,mul954,s924);   adder a954(s924,mul955,s925);   adder a955(s925,mul956,s926);   adder a956(s926,mul957,s927);   adder a957(s927,mul958,s928);   adder a958(s928,mul959,s929);   
	adder a960(mul960,mul961,s930);   adder a961(s930,mul962,s931);   adder a962(s931,mul963,s932);   adder a963(s932,mul964,s933);   adder a964(s933,mul965,s934);   adder a965(s934,mul966,s935);   adder a966(s935,mul967,s936);   adder a967(s936,mul968,s937);   adder a968(s937,mul969,s938);   adder a969(s938,mul970,s939);   adder a970(s939,mul971,s940);   adder a971(s940,mul972,s941);   adder a972(s941,mul973,s942);   adder a973(s942,mul974,s943);   adder a974(s943,mul975,s944);   adder a975(s944,mul976,s945);   adder a976(s945,mul977,s946);   adder a977(s946,mul978,s947);   adder a978(s947,mul979,s948);   adder a979(s948,mul980,s949);   adder a980(s949,mul981,s950);   adder a981(s950,mul982,s951);   adder a982(s951,mul983,s952);   adder a983(s952,mul984,s953);   adder a984(s953,mul985,s954);   adder a985(s954,mul986,s955);   adder a986(s955,mul987,s956);   adder a987(s956,mul988,s957);   adder a988(s957,mul989,s958);   adder a989(s958,mul990,s959);   adder a990(s959,mul991,s960);   
	adder a992(mul992,mul993,s961);   adder a993(s961,mul994,s962);   adder a994(s962,mul995,s963);   adder a995(s963,mul996,s964);   adder a996(s964,mul997,s965);   adder a997(s965,mul998,s966);   adder a998(s966,mul999,s967);   adder a999(s967,mul1000,s968);   adder a1000(s968,mul1001,s969);   adder a1001(s969,mul1002,s970);   adder a1002(s970,mul1003,s971);   adder a1003(s971,mul1004,s972);   adder a1004(s972,mul1005,s973);   adder a1005(s973,mul1006,s974);   adder a1006(s974,mul1007,s975);   adder a1007(s975,mul1008,s976);   adder a1008(s976,mul1009,s977);   adder a1009(s977,mul1010,s978);   adder a1010(s978,mul1011,s979);   adder a1011(s979,mul1012,s980);   adder a1012(s980,mul1013,s981);   adder a1013(s981,mul1014,s982);   adder a1014(s982,mul1015,s983);   adder a1015(s983,mul1016,s984);   adder a1016(s984,mul1017,s985);   adder a1017(s985,mul1018,s986);   adder a1018(s986,mul1019,s987);   adder a1019(s987,mul1020,s988);   adder a1020(s988,mul1021,s989);   adder a1021(s989,mul1022,s990);   adder a1022(s990,mul1023,s991);  
	
	assign address = address_reg + 5'b00001;
	
	always@(posedge clk)
		begin
			if(reset == 1'b1)
				begin
					loaded_flag <= 1'b0;
					address_reg <= 5'b11111;
				end
			else if(loaded_flag == 1'b0)
				begin
						for(i = 0;i < 32; i = i + 1)
							begin
								A[index_A][i] <= A_wire[1023 - 10'd32*i -: 10'd32];
								B[index_B][i] <= B_wire[1023 - 10'd32*i -: 10'd32];
							end
						if(index_A == 5'b11111)
							begin
								loaded_flag = 1'b1;
							end
				end
			else
				begin
					C[address][0] <= s30;
					C[address][1] <= s61;
					C[address][2] <= s92;
					C[address][3] <= sum3;
					C[address][4] <= sum4;
					C[address][5] <= sum5;
					C[address][6] <= sum6;
					C[address][7] <= sum7;
					C[address][8] <= sum8;
					C[address][9] <= sum9;
					C[address][10] <= sum10;
					C[address][11] <= sum11;
					C[address][12] <= sum12;
					C[address][13] <= sum13;
					C[address][14] <= sum14;
					C[address][15] <= sum15;
					C[address][16] <= sum16;
					C[address][17] <= sum17;
					C[address][18] <= sum18;
					C[address][19] <= sum19;
					C[address][20] <= sum20;
					C[address][21] <= sum21;
					C[address][22] <= sum22;
					C[address][23] <= sum23;
					C[address][24] <= sum24;
					C[address][25] <= sum25;
					C[address][26] <= sum26;
					C[address][27] <= sum27;
					C[address][28] <= sum28;
					C[address][29] <= sum29;
					C[address][30] <= sum30;
					C[address][31] <= sum31;
					*/
					for(i = 0; i < 32; i = i + 1)
						begin
							out[1023 - 10'd32*i -: 10'd32] <= C[address][i];
							$display("out: %d", out[1023 - 10'd32*i -: 10'd32]);
						end
//					write_out <= 1'b1;
					address_reg <= address;					
					out_address <= address;
					select_line_out <= select_line_in;
				end
		end
endmodule

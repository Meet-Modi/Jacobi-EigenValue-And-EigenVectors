`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   01:22:53 11/14/2018
// Design Name:   Matrix_Multiply_32
// Module Name:   C:/MEET/PROJECTS/COLASS/Final_32/Matrix_Multiply_32_tb.v
// Project Name:  Final_32
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Matrix_Multiply_32
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Matrix_Multiply_32_tb;

	// Inputs
	reg select_line_in;
	reg [1023:0] A_wire;
	reg [1023:0] B_wire;
	reg [4:0] index_A;
	reg [4:0] index_B;
	reg clk;
	reg reset;

	// Outputs
	wire [1023:0] out;
	wire [4:0] out_address;
	wire select_line_out;
	wire write_data;

	// Instantiate the Unit Under Test (UUT)
	Matrix_Multiply_32 uut (
		.select_line_in(select_line_in), 
		.A_wire(A_wire), 
		.B_wire(B_wire), 
		.index_A(index_A), 
		.index_B(index_B), 
		.clk(clk), 
		.reset(reset), 
		.out(out), 
		.out_address(out_address), 
		.select_line_out(select_line_out), 
		.write_data(write_data)
	);

	initial begin
		select_line_in = 0;
		A_wire = 0;
		B_wire = 0;
		index_A = 0;
		index_B = 0;
		clk = 0;
		reset = 0;
		
		#3 reset = 1'b1;
		#3 reset = 1'b0;
	
		A_wire = 1024'b0000000000000000000000000001000000000000000000000000000001111000000000000000000000000000100010110000000000000000000000001000011100000000000000000000000011101010000000000000000000000000111011000000000000000000000000001010110100000000000000000000000001000111000000000000000000000000011111100000000000000000000000001000001000000000000000000000000000100001000000000000000000000000111100010000000000000000000000000010100000000000000000000000000001001010000000000000000000000000111110100000000000000000000000000100110000000000000000000000000001100010000000000000000000000000001110100000000000000000000000000101111100000000000000000000000001111101000000000000000000000000111001010000000000000000000000000010000100000000000000000000000000100001000000000000000000000000110101010000000000000000000000001010001100000000000000000000000000000011000000000000000000000000111011100000000000000000000000001111001000000000000000000000000001110001000000000000000000000000000110000000000000000000000000000100011100000000000000000000000001101110;
		B_wire = 1024'b0000000000000000000000000001000000000000000000000000000001111000000000000000000000000000100010110000000000000000000000001000011100000000000000000000000011101010000000000000000000000000111011000000000000000000000000001010110100000000000000000000000001000111000000000000000000000000011111100000000000000000000000001000001000000000000000000000000000100001000000000000000000000000111100010000000000000000000000000010100000000000000000000000000001001010000000000000000000000000111110100000000000000000000000000100110000000000000000000000000001100010000000000000000000000000001110100000000000000000000000000101111100000000000000000000000001111101000000000000000000000000111001010000000000000000000000000010000100000000000000000000000000100001000000000000000000000000110101010000000000000000000000001010001100000000000000000000000000000011000000000000000000000000111011100000000000000000000000001111001000000000000000000000000001110001000000000000000000000000000110000000000000000000000000000100011100000000000000000000000001101110;
		
		index_A = 5'd0;
		index_B = 5'd0;

		#10
    	index_A = 5'd1;
		index_B = 5'd1;

		#10

		index_A = 5'd2;
		index_B = 5'd2;
		
		#10
    		
		index_A = 5'd3;
		index_B = 5'd3;

		#10
		
		index_A = 5'd4;
		index_B = 5'd4;

		#10
		
		index_A = 5'd5;
		index_B = 5'd5;

		#10
		
		index_A = 5'd6;
		index_B = 5'd6;

		#10
		
		index_A = 5'd7;
		index_B = 5'd7;
		
		#10
		
		index_A = 5'd8;
		index_B = 5'd8;
		
		#10
		
		index_A = 5'd9;
		index_B = 5'd9;
		
		#10
		
		index_A = 5'd10;
		index_B = 5'd10;


		#10
		
		index_A = 5'd11;
		index_B = 5'd11;
		
		#10
		
		index_A = 5'd12;
		index_B = 5'd12;

		#10
		
		index_A = 5'd13;
		index_B = 5'd13;
		
		#10
		
		index_A = 5'd14;
		index_B = 5'd14;

		#10
		
		index_A = 5'd15;
		index_B = 5'd15;

		#10
		
		index_A = 5'd16;
		index_B = 5'd16;

		#10
		
		index_A = 5'd17;
		index_B = 5'd17;

		#10
		
		index_A = 5'd18;
		index_B = 5'd18;

		#10
		
		index_A = 5'd19;
		index_B = 5'd19;

		#10
		
		index_A = 5'd20;
		index_B = 5'd20;

		#10
		
		index_A = 5'd21;
		index_B = 5'd21;

		#10
		
		index_A = 5'd22;
		index_B = 5'd22;

		#10
		
		index_A = 5'd23;
		index_B = 5'd23;

		#10
		
		index_A = 5'd24;
		index_B = 5'd24;

		#10
		
		index_A = 5'd25;
		index_B = 5'd25;

		#10
		
		index_A = 5'd26;
		index_B = 5'd26;

		#10
		
		index_A = 5'd27;
		index_B = 5'd27;

		#10
		
		index_A = 5'd28;
		index_B = 5'd28;

		#10
		
		index_A = 5'd29;
		index_B = 5'd29;

		#10
		
		index_A = 5'd30;
		index_B = 5'd30;

		#10
		
		index_A = 5'd31;
		index_B = 5'd31;

	end
      always #5 clk = ~clk;

endmodule


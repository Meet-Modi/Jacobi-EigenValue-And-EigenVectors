`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   01:32:21 11/14/2018
// Design Name:   RAM
// Module Name:   C:/MEET/PROJECTS/COLASS/Final_32/RAM_tb.v
// Project Name:  Final_32
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: RAM
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module RAM_tb;

	// Inputs
	reg clk;
	reg reset;
	reg ena;
	reg read_write;
	reg [4:0] address_1;
	reg [4:0] address_2;
	reg [1023:0] data_in_1;
	reg [1023:0] data_in_2;
	reg data_in_mux;
	reg data_out_mux;
	reg address_mux;

	// Outputs
	wire [1023:0] data_out_1;
	wire [1023:0] data_out_2;

	// Instantiate the Unit Under Test (UUT)
	RAM uut (
		.clk(clk), 
		.reset(reset), 
		.ena(ena), 
		.read_write(read_write), 
		.address_1(address_1), 
		.address_2(address_2), 
		.data_in_1(data_in_1), 
		.data_in_2(data_in_2), 
		.data_out_1(data_out_1), 
		.data_out_2(data_out_2), 
		.data_in_mux(data_in_mux), 
		.data_out_mux(data_out_mux), 
		.address_mux(address_mux)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1'b0;
		
		ena = 1'b1;
		read_write = 1'b1;
		address_1 = 5'd0;
		address_2 = 5'd0;
		data_in_1 = 1024'b0000000000000000000000000001000000000000000000000000000001111000000000000000000000000000100010110000000000000000000000001000011100000000000000000000000011101010000000000000000000000000111011000000000000000000000000001010110100000000000000000000000001000111000000000000000000000000011111100000000000000000000000001000001000000000000000000000000000100001000000000000000000000000111100010000000000000000000000000010100000000000000000000000000001001010000000000000000000000000111110100000000000000000000000000100110000000000000000000000000001100010000000000000000000000000001110100000000000000000000000000101111100000000000000000000000001111101000000000000000000000000111001010000000000000000000000000010000100000000000000000000000000100001000000000000000000000000110101010000000000000000000000001010001100000000000000000000000000000011000000000000000000000000111011100000000000000000000000001111001000000000000000000000000001110001000000000000000000000000000110000000000000000000000000000100011100000000000000000000000001101110;
		data_in_2 = 1024'b1000000000000000000000000000100000000000000000000000000000111100000000000000000000000000010001011000000000000000000000000100001110000000000000000000000001110101000000000000000000000000011101100000000000000000000000000101011010000000000000000000000000100011100000000000000000000000001111110000000000000000000000000100000100000000000000000000000000010000100000000000000000000000011110001000000000000000000000000001010000000000000000000000000000100101000000000000000000000000011111010000000000000000000000000010011000000000000000000000000000110001000000000000000000000000000111010000000000000000000000000010111110000000000000000000000000111110100000000000000000000000011100101000000000000000000000000001000010000000000000000000000000010000100000000000000000000000011010101000000000000000000000000101000110000000000000000000000000000001100000000000000000000000011101110000000000000000000000000111100100000000000000000000000000111000100000000000000000000000000011000000000000000000000000000010001110000000000000000000000000110111;;
		data_in_mux = 1'b0;
		data_out_mux = 1'b0;
		address_mux = 1'b0;
		
		#15
		ena = 1'b1;
		reset = 1'b1;
		read_write = 1'b1;
		address_1 = 5'd0;
		address_2 = 5'd0;
		data_in_mux = 1'b1;
		data_out_mux = 1'b0;
		address_mux = 1'b1;	
		
		
		#15
		ena = 1'b1;
		reset = 1'b1;
		read_write = 1'b0;
		address_1 = 5'd0;
		address_2 = 5'd0;
		data_in_mux = 1'b0;
		data_out_mux = 1'b0;
		address_mux = 1'b0;	
		
		#15
		ena = 1'b1;
		reset = 1'b1;
		read_write = 1'b0;
		address_1 = 5'd0;
		address_2 = 5'd0;
		data_in_mux = 1'b1;
		data_out_mux = 1'b1;
		address_mux = 1'b1;	
		
		
	end
      always #5 clk = ~clk;
endmodule


`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   00:58:53 11/13/2018
// Design Name:   Matrix_Multiply_32_final
// Module Name:   C:/MEET/PROJECTS/COLASS/Final_32/Matrix_Multiply_32_final_tb.v
// Project Name:  Final_32
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Matrix_Multiply_32_final
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Matrix_Multiply_32_final_tb;

	// Inputs
	reg [1023:0] A_wire;
	reg [1023:0] B_wire;
	reg clk;
	reg reset;
	reg [4:0] index_A;
	reg [4:0] index_B;

	// Outputs
	wire [1023:0] Answer;

	// Instantiate the Unit Under Test (UUT)
	Matrix_Multiply_32_final uut (
		.Answer(Answer), 
		.A_wire(A_wire), 
		.B_wire(B_wire), 
		.clk(clk), 
		.reset(reset), 
		.index_A(index_A), 
		.index_B(index_B)
	);

		initial begin
		// Initialize Inputs
		A_wire = 0;
		B_wire = 0;
		clk = 0;
		reset = 0;
		index_A = 5'd0;
		index_B = 5'd0;
		
		#3 reset = 1'b1;
		#3 reset = 1'b0;
		
		/*A_wire = 1024'b0;
		B_wire = 1024'b0;
		*/
		
		A_wire = 1024'b000000000000000000000000000010000000000000000000000000000011110000000000000000000000000001000101100000000000000000000000010000111000000000000000000000000111010100000000000000000000000001110110000000000000000000000000010101101000000000000000000000000010001110000000000000000000000000111111000000000000000000000000010000010000000000000000000000000001000010000000000000000000000001111000100000000000000000000000000101000000000000000000000000000010010100000000000000000000000001111101000000000000000000000000001001100000000000000000000000000011000100000000000000000000000000011101000000000000000000000000001011111000000000000000000000000011111010000000000000000000000001110010100000000000000000000000000100001000000000000000000000000001000010000000000000000000000001101010100000000000000000000000010100011000000000000000000000000000000110000000000000000000000001110111000000000000000000000000011110010000000000000000000000000011100010000000000000000000000000001100000000000000000000000000001000111000000000000000000000000011011;
		B_wire = 1024'b000000000000000000000000000010000000000000000000000000000011110000000000000000000000000001000101100000000000000000000000010000111000000000000000000000000111010100000000000000000000000001110110000000000000000000000000010101101000000000000000000000000010001110000000000000000000000000111111000000000000000000000000010000010000000000000000000000000001000010000000000000000000000001111000100000000000000000000000000101000000000000000000000000000010010100000000000000000000000001111101000000000000000000000000001001100000000000000000000000000011000100000000000000000000000000011101000000000000000000000000001011111000000000000000000000000011111010000000000000000000000001110010100000000000000000000000000100001000000000000000000000000001000010000000000000000000000001101010100000000000000000000000010100011000000000000000000000000000000110000000000000000000000001110111000000000000000000000000011110010000000000000000000000000011100010000000000000000000000000001100000000000000000000000000001000111000000000000000000000000011011;
		index_A = 5'd0;
		index_B = 5'd0;

		#10
    	index_A = 5'd1;
		index_B = 5'd1;

		#10

		index_A = 5'd2;
		index_B = 5'd2;
		
		#10
    		
		index_A = 5'd3;
		index_B = 5'd3;

		#10
		
		index_A = 5'd4;
		index_B = 5'd4;

		#10
		
		index_A = 5'd5;
		index_B = 5'd5;

		#10
		
		index_A = 5'd6;
		index_B = 5'd6;

		#10
		
		index_A = 5'd7;
		index_B = 5'd7;
		
		#10
		
		index_A = 5'd8;
		index_B = 5'd8;
		
		#10
		
		index_A = 5'd9;
		index_B = 5'd9;

		#10
		
		index_A = 5'd11;
		index_B = 5'd11;
		
		#10
		
		index_A = 5'd12;
		index_B = 5'd12;

		#10
		
		index_A = 5'd13;
		index_B = 5'd13;
		
		#10
		
		index_A = 5'd14;
		index_B = 5'd14;

		#10
		
		index_A = 5'd15;
		index_B = 5'd15;

		#10
		
		index_A = 5'd16;
		index_B = 5'd16;

		#10
		
		index_A = 5'd17;
		index_B = 5'd17;

		#10
		
		index_A = 5'd18;
		index_B = 5'd18;

		#10
		
		index_A = 5'd19;
		index_B = 5'd19;

		#10
		
		index_A = 5'd20;
		index_B = 5'd20;

		#10
		
		index_A = 5'd21;
		index_B = 5'd21;

		#10
		
		index_A = 5'd22;
		index_B = 5'd22;

		#10
		
		index_A = 5'd23;
		index_B = 5'd23;

		#10
		
		index_A = 5'd24;
		index_B = 5'd24;

		#10
		
		index_A = 5'd25;
		index_B = 5'd25;

		#10
		
		index_A = 5'd26;
		index_B = 5'd26;

		#10
		
		index_A = 5'd27;
		index_B = 5'd27;

		#10
		
		index_A = 5'd28;
		index_B = 5'd28;

		#10
		
		index_A = 5'd29;
		index_B = 5'd29;

		#10
		
		index_A = 5'd30;
		index_B = 5'd30;

		#10
		
		index_A = 5'd31;
		index_B = 5'd31;

	end
      always #5 clk = ~clk;
endmodule



